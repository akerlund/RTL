////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2021 Fredrik Åkerlund
// https://github.com/akerlund/RTL
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <https://www.gnu.org/licenses/>.
//
// Description:
//
////////////////////////////////////////////////////////////////////////////////

`default_nettype none

module gray_to_bin #(
    parameter WIDTH_P = -1
  )(
    input  wire  [WIDTH_P-1 : 0] gray,
    output logic [WIDTH_P-1 : 0] bin
  );

  genvar i;

  generate
    for (i = 0; i < WIDTH_P; i++) begin
      assign bin[i] = ^gray[WIDTH_P-1 : i];
    end
  endgenerate

endmodule

`default_nettype wire
