package gf_ref_pkg;

localparam int M_C        = 256;
localparam int REF_SIZE_C = 16;

localparam logic [M_C-1 : 0] GF_ADD_C [REF_SIZE_C] [3] = '{
  '{91,198,157},
  '{217,121,160},
  '{233,204,37},
  '{222,16,206},
  '{249,88,161},
  '{88,104,48},
  '{202,228,46},
  '{85,228,177},
  '{98,85,55},
  '{105,25,112},
  '{243,250,9},
  '{49,198,247},
  '{246,111,153},
  '{206,107,165},
  '{127,174,209},
  '{199,83,148}
};

localparam logic [M_C-1 : 0] GF_MUL_C [REF_SIZE_C] [3] = '{
  '{2,185,105},
  '{144,160,223},
  '{51,148,57},
  '{103,24,63},
  '{130,186,241},
  '{152,218,253},
  '{97,21,180},
  '{243,9,42},
  '{205,205,96},
  '{150,66,141},
  '{201,191,12},
  '{16,182,149},
  '{148,55,95},
  '{195,89,35},
  '{70,112,36},
  '{217,185,233}
};

localparam logic [M_C-1 : 0] GF_DIV_C [REF_SIZE_C] [3] = '{
  '{110,63,145},
  '{102,188,145},
  '{166,11,145},
  '{206,78,145},
  '{57,38,145},
  '{158,86,145},
  '{116,79,145},
  '{215,174,145},
  '{35,109,145},
  '{162,108,145},
  '{102,1,145},
  '{42,104,145},
  '{85,140,145},
  '{129,225,145},
  '{160,175,145},
  '{97,96,145}
};

endpackage
