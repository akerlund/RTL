`include "vip_axi4s_if.sv"
`include "vip_axi4s_pkg.sv"
