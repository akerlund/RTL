`include "uvm_macros.svh"
import uvm_pkg::*;

`include "axi4s_m2s_2m_arbiter.sv"
