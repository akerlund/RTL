////////////////////////////////////////////////////////////////////////////////
//
// Copyright 2020 Fredrik Åkerlund
//
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either
// version 2.1 of the License, or (at your option) any later version.
//
// This library is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public
// License along with this library; if not, write to the Free Software
// Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA 02110-1301, USA
//
// Description:
//
////////////////////////////////////////////////////////////////////////////////

`ifndef CORDIC_TEST_ANGLES_PKG
`define CORDIC_TEST_ANGLES_PKG

package cordic_test_angles_pkg;

  logic [31 : 0] test_angles [360] = {
    32'b00000000000000000000000000000000,
    32'b00000000101101100000101101100001,
    32'b00000001011011000001011011000001,
    32'b00000010001000100010001000100010,
    32'b00000010110110000010110110000011,
    32'b00000011100011100011100011100100,
    32'b00000100010001000100010001000100,
    32'b00000100111110100100111110100101,
    32'b00000101101100000101101100000110,
    32'b00000110011001100110011001100110,
    32'b00000111000111000111000111000111,
    32'b00000111110100100111110100101000,
    32'b00001000100010001000100010001001,
    32'b00001001001111101001001111101001,
    32'b00001001111101001001111101001010,
    32'b00001010101010101010101010101011,
    32'b00001011011000001011011000001011,
    32'b00001100000101101100000101101100,
    32'b00001100110011001100110011001101,
    32'b00001101100000101101100000101110,
    32'b00001110001110001110001110001110,
    32'b00001110111011101110111011101111,
    32'b00001111101001001111101001010000,
    32'b00010000010110110000010110110000,
    32'b00010001000100010001000100010001,
    32'b00010001110001110001110001110010,
    32'b00010010011111010010011111010010,
    32'b00010011001100110011001100110011,
    32'b00010011111010010011111010010100,
    32'b00010100100111110100100111110101,
    32'b00010101010101010101010101010101,
    32'b00010110000010110110000010110110,
    32'b00010110110000010110110000010111,
    32'b00010111011101110111011101110111,
    32'b00011000001011011000001011011000,
    32'b00011000111000111000111000111001,
    32'b00011001100110011001100110011010,
    32'b00011010010011111010010011111010,
    32'b00011011000001011011000001011011,
    32'b00011011101110111011101110111100,
    32'b00011100011100011100011100011100,
    32'b00011101001001111101001001111101,
    32'b00011101110111011101110111011110,
    32'b00011110100100111110100100111111,
    32'b00011111010010011111010010011111,
    32'b00100000000000000000000000000000,
    32'b00100000101101100000101101100001,
    32'b00100001011011000001011011000001,
    32'b00100010001000100010001000100010,
    32'b00100010110110000010110110000011,
    32'b00100011100011100011100011100100,
    32'b00100100010001000100010001000100,
    32'b00100100111110100100111110100101,
    32'b00100101101100000101101100000110,
    32'b00100110011001100110011001100110,
    32'b00100111000111000111000111000111,
    32'b00100111110100100111110100101000,
    32'b00101000100010001000100010001001,
    32'b00101001001111101001001111101001,
    32'b00101001111101001001111101001010,
    32'b00101010101010101010101010101011,
    32'b00101011011000001011011000001011,
    32'b00101100000101101100000101101100,
    32'b00101100110011001100110011001101,
    32'b00101101100000101101100000101110,
    32'b00101110001110001110001110001110,
    32'b00101110111011101110111011101111,
    32'b00101111101001001111101001010000,
    32'b00110000010110110000010110110000,
    32'b00110001000100010001000100010001,
    32'b00110001110001110001110001110010,
    32'b00110010011111010010011111010010,
    32'b00110011001100110011001100110011,
    32'b00110011111010010011111010010100,
    32'b00110100100111110100100111110101,
    32'b00110101010101010101010101010101,
    32'b00110110000010110110000010110110,
    32'b00110110110000010110110000010111,
    32'b00110111011101110111011101110111,
    32'b00111000001011011000001011011000,
    32'b00111000111000111000111000111001,
    32'b00111001100110011001100110011010,
    32'b00111010010011111010010011111010,
    32'b00111011000001011011000001011011,
    32'b00111011101110111011101110111100,
    32'b00111100011100011100011100011100,
    32'b00111101001001111101001001111101,
    32'b00111101110111011101110111011110,
    32'b00111110100100111110100100111111,
    32'b00111111010010011111010010011111,
    32'b01000000000000000000000000000000,
    32'b01000000101101100000101101100001,
    32'b01000001011011000001011011000001,
    32'b01000010001000100010001000100010,
    32'b01000010110110000010110110000011,
    32'b01000011100011100011100011100100,
    32'b01000100010001000100010001000100,
    32'b01000100111110100100111110100101,
    32'b01000101101100000101101100000110,
    32'b01000110011001100110011001100110,
    32'b01000111000111000111000111000111,
    32'b01000111110100100111110100101000,
    32'b01001000100010001000100010001001,
    32'b01001001001111101001001111101001,
    32'b01001001111101001001111101001010,
    32'b01001010101010101010101010101011,
    32'b01001011011000001011011000001011,
    32'b01001100000101101100000101101100,
    32'b01001100110011001100110011001101,
    32'b01001101100000101101100000101110,
    32'b01001110001110001110001110001110,
    32'b01001110111011101110111011101111,
    32'b01001111101001001111101001010000,
    32'b01010000010110110000010110110000,
    32'b01010001000100010001000100010001,
    32'b01010001110001110001110001110010,
    32'b01010010011111010010011111010010,
    32'b01010011001100110011001100110011,
    32'b01010011111010010011111010010100,
    32'b01010100100111110100100111110101,
    32'b01010101010101010101010101010101,
    32'b01010110000010110110000010110110,
    32'b01010110110000010110110000010111,
    32'b01010111011101110111011101110111,
    32'b01011000001011011000001011011000,
    32'b01011000111000111000111000111001,
    32'b01011001100110011001100110011010,
    32'b01011010010011111010010011111010,
    32'b01011011000001011011000001011011,
    32'b01011011101110111011101110111100,
    32'b01011100011100011100011100011100,
    32'b01011101001001111101001001111101,
    32'b01011101110111011101110111011110,
    32'b01011110100100111110100100111111,
    32'b01011111010010011111010010011111,
    32'b01100000000000000000000000000000,
    32'b01100000101101100000101101100001,
    32'b01100001011011000001011011000001,
    32'b01100010001000100010001000100010,
    32'b01100010110110000010110110000011,
    32'b01100011100011100011100011100100,
    32'b01100100010001000100010001000100,
    32'b01100100111110100100111110100101,
    32'b01100101101100000101101100000110,
    32'b01100110011001100110011001100110,
    32'b01100111000111000111000111000111,
    32'b01100111110100100111110100101000,
    32'b01101000100010001000100010001001,
    32'b01101001001111101001001111101001,
    32'b01101001111101001001111101001010,
    32'b01101010101010101010101010101011,
    32'b01101011011000001011011000001011,
    32'b01101100000101101100000101101100,
    32'b01101100110011001100110011001101,
    32'b01101101100000101101100000101110,
    32'b01101110001110001110001110001110,
    32'b01101110111011101110111011101111,
    32'b01101111101001001111101001010000,
    32'b01110000010110110000010110110000,
    32'b01110001000100010001000100010001,
    32'b01110001110001110001110001110010,
    32'b01110010011111010010011111010010,
    32'b01110011001100110011001100110011,
    32'b01110011111010010011111010010100,
    32'b01110100100111110100100111110101,
    32'b01110101010101010101010101010101,
    32'b01110110000010110110000010110110,
    32'b01110110110000010110110000010111,
    32'b01110111011101110111011101110111,
    32'b01111000001011011000001011011000,
    32'b01111000111000111000111000111001,
    32'b01111001100110011001100110011010,
    32'b01111010010011111010010011111010,
    32'b01111011000001011011000001011011,
    32'b01111011101110111011101110111100,
    32'b01111100011100011100011100011100,
    32'b01111101001001111101001001111101,
    32'b01111101110111011101110111011110,
    32'b01111110100100111110100100111111,
    32'b01111111010010011111010010011111,
    32'b10000000000000000000000000000000,
    32'b10000000101101100000101101100001,
    32'b10000001011011000001011011000001,
    32'b10000010001000100010001000100010,
    32'b10000010110110000010110110000011,
    32'b10000011100011100011100011100100,
    32'b10000100010001000100010001000100,
    32'b10000100111110100100111110100101,
    32'b10000101101100000101101100000110,
    32'b10000110011001100110011001100110,
    32'b10000111000111000111000111000111,
    32'b10000111110100100111110100101000,
    32'b10001000100010001000100010001001,
    32'b10001001001111101001001111101001,
    32'b10001001111101001001111101001010,
    32'b10001010101010101010101010101011,
    32'b10001011011000001011011000001011,
    32'b10001100000101101100000101101100,
    32'b10001100110011001100110011001101,
    32'b10001101100000101101100000101110,
    32'b10001110001110001110001110001110,
    32'b10001110111011101110111011101111,
    32'b10001111101001001111101001010000,
    32'b10010000010110110000010110110000,
    32'b10010001000100010001000100010001,
    32'b10010001110001110001110001110010,
    32'b10010010011111010010011111010010,
    32'b10010011001100110011001100110011,
    32'b10010011111010010011111010010100,
    32'b10010100100111110100100111110101,
    32'b10010101010101010101010101010101,
    32'b10010110000010110110000010110110,
    32'b10010110110000010110110000010111,
    32'b10010111011101110111011101110111,
    32'b10011000001011011000001011011000,
    32'b10011000111000111000111000111001,
    32'b10011001100110011001100110011010,
    32'b10011010010011111010010011111010,
    32'b10011011000001011011000001011011,
    32'b10011011101110111011101110111100,
    32'b10011100011100011100011100011100,
    32'b10011101001001111101001001111101,
    32'b10011101110111011101110111011110,
    32'b10011110100100111110100100111111,
    32'b10011111010010011111010010011111,
    32'b10100000000000000000000000000000,
    32'b10100000101101100000101101100001,
    32'b10100001011011000001011011000001,
    32'b10100010001000100010001000100010,
    32'b10100010110110000010110110000011,
    32'b10100011100011100011100011100100,
    32'b10100100010001000100010001000100,
    32'b10100100111110100100111110100101,
    32'b10100101101100000101101100000110,
    32'b10100110011001100110011001100110,
    32'b10100111000111000111000111000111,
    32'b10100111110100100111110100101000,
    32'b10101000100010001000100010001001,
    32'b10101001001111101001001111101001,
    32'b10101001111101001001111101001010,
    32'b10101010101010101010101010101011,
    32'b10101011011000001011011000001011,
    32'b10101100000101101100000101101100,
    32'b10101100110011001100110011001101,
    32'b10101101100000101101100000101110,
    32'b10101110001110001110001110001110,
    32'b10101110111011101110111011101111,
    32'b10101111101001001111101001010000,
    32'b10110000010110110000010110110000,
    32'b10110001000100010001000100010001,
    32'b10110001110001110001110001110010,
    32'b10110010011111010010011111010010,
    32'b10110011001100110011001100110011,
    32'b10110011111010010011111010010100,
    32'b10110100100111110100100111110101,
    32'b10110101010101010101010101010101,
    32'b10110110000010110110000010110110,
    32'b10110110110000010110110000010111,
    32'b10110111011101110111011101110111,
    32'b10111000001011011000001011011000,
    32'b10111000111000111000111000111001,
    32'b10111001100110011001100110011010,
    32'b10111010010011111010010011111010,
    32'b10111011000001011011000001011011,
    32'b10111011101110111011101110111100,
    32'b10111100011100011100011100011100,
    32'b10111101001001111101001001111101,
    32'b10111101110111011101110111011110,
    32'b10111110100100111110100100111111,
    32'b10111111010010011111010010011111,
    32'b11000000000000000000000000000000,
    32'b11000000101101100000101101100001,
    32'b11000001011011000001011011000001,
    32'b11000010001000100010001000100010,
    32'b11000010110110000010110110000011,
    32'b11000011100011100011100011100100,
    32'b11000100010001000100010001000100,
    32'b11000100111110100100111110100101,
    32'b11000101101100000101101100000110,
    32'b11000110011001100110011001100110,
    32'b11000111000111000111000111000111,
    32'b11000111110100100111110100101000,
    32'b11001000100010001000100010001001,
    32'b11001001001111101001001111101001,
    32'b11001001111101001001111101001010,
    32'b11001010101010101010101010101011,
    32'b11001011011000001011011000001011,
    32'b11001100000101101100000101101100,
    32'b11001100110011001100110011001101,
    32'b11001101100000101101100000101110,
    32'b11001110001110001110001110001110,
    32'b11001110111011101110111011101111,
    32'b11001111101001001111101001010000,
    32'b11010000010110110000010110110000,
    32'b11010001000100010001000100010001,
    32'b11010001110001110001110001110010,
    32'b11010010011111010010011111010010,
    32'b11010011001100110011001100110011,
    32'b11010011111010010011111010010100,
    32'b11010100100111110100100111110101,
    32'b11010101010101010101010101010101,
    32'b11010110000010110110000010110110,
    32'b11010110110000010110110000010111,
    32'b11010111011101110111011101110111,
    32'b11011000001011011000001011011000,
    32'b11011000111000111000111000111001,
    32'b11011001100110011001100110011010,
    32'b11011010010011111010010011111010,
    32'b11011011000001011011000001011011,
    32'b11011011101110111011101110111100,
    32'b11011100011100011100011100011100,
    32'b11011101001001111101001001111101,
    32'b11011101110111011101110111011110,
    32'b11011110100100111110100100111111,
    32'b11011111010010011111010010011111,
    32'b11100000000000000000000000000000,
    32'b11100000101101100000101101100001,
    32'b11100001011011000001011011000001,
    32'b11100010001000100010001000100010,
    32'b11100010110110000010110110000011,
    32'b11100011100011100011100011100100,
    32'b11100100010001000100010001000100,
    32'b11100100111110100100111110100101,
    32'b11100101101100000101101100000110,
    32'b11100110011001100110011001100110,
    32'b11100111000111000111000111000111,
    32'b11100111110100100111110100101000,
    32'b11101000100010001000100010001001,
    32'b11101001001111101001001111101001,
    32'b11101001111101001001111101001010,
    32'b11101010101010101010101010101011,
    32'b11101011011000001011011000001011,
    32'b11101100000101101100000101101100,
    32'b11101100110011001100110011001101,
    32'b11101101100000101101100000101110,
    32'b11101110001110001110001110001110,
    32'b11101110111011101110111011101111,
    32'b11101111101001001111101001010000,
    32'b11110000010110110000010110110000,
    32'b11110001000100010001000100010001,
    32'b11110001110001110001110001110010,
    32'b11110010011111010010011111010010,
    32'b11110011001100110011001100110011,
    32'b11110011111010010011111010010100,
    32'b11110100100111110100100111110101,
    32'b11110101010101010101010101010101,
    32'b11110110000010110110000010110110,
    32'b11110110110000010110110000010111,
    32'b11110111011101110111011101110111,
    32'b11111000001011011000001011011000,
    32'b11111000111000111000111000111001,
    32'b11111001100110011001100110011010,
    32'b11111010010011111010010011111010,
    32'b11111011000001011011000001011011,
    32'b11111011101110111011101110111100,
    32'b11111100011100011100011100011100,
    32'b11111101001001111101001001111101,
    32'b11111101110111011101110111011110,
    32'b11111110100100111110100100111111,
    32'b11111111010010011111010010011111
  };

endpackage

`endif
