////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2020 Fredrik Åkerlund
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <https://www.gnu.org/licenses/>.
//
// Description:
//
////////////////////////////////////////////////////////////////////////////////

// There is a gain of 3 bits, therefore:
// Maximum input size is 63.984375
// Minimum input size is -64.0
// Maximum output size is 511.984375
// Minimum output size is -512.0
//
// Smallest output is -171.421875
// Largest  output is 171.421875

package tb_fft_N8_Q10_6_test_data_pkg;

localparam int nr_of_tests_c   = 64;
localparam int data_width_c    = 16;
localparam int nr_of_samples_c = 8;
localparam int nr_of_n_bits_c  = 10;
localparam int nr_of_q_bits_c  = 6;

logic [15 : 0] x_test_data_re [nr_of_tests_c][8] = {
  // x_re_0 = [-38.390625, -36.203125, 22.296875, 36.59375, 5.640625, -5.28125, 22.625, -44.0]
  {
    16'b1111011001100111,  // -38.390625
    16'b1111011011110011,  // -36.203125
    16'b0000010110010011,  // 22.296875
    16'b0000100100100110,  // 36.59375
    16'b0000000101101001,  // 5.640625
    16'b1111111010101110,  // -5.28125
    16'b0000010110101000,  // 22.625
    16'b1111010100000000   // -44.0
  },
  // x_re_1 = [-21.609375, 30.390625, 35.453125, -12.140625, 52.953125, -36.546875, 59.96875, -2.78125]
  {
    16'b1111101010011001,  // -21.609375
    16'b0000011110011001,  // 30.390625
    16'b0000100011011101,  // 35.453125
    16'b1111110011110111,  // -12.140625
    16'b0000110100111101,  // 52.953125
    16'b1111011011011101,  // -36.546875
    16'b0000111011111110,  // 59.96875
    16'b1111111101001110   // -2.78125
  },
  // x_re_2 = [36.578125, 56.828125, -52.875, -41.453125, -16.296875, 48.59375, -8.65625, 51.09375]
  {
    16'b0000100100100101,  // 36.578125
    16'b0000111000110101,  // 56.828125
    16'b1111001011001000,  // -52.875
    16'b1111010110100011,  // -41.453125
    16'b1111101111101101,  // -16.296875
    16'b0000110000100110,  // 48.59375
    16'b1111110111010110,  // -8.65625
    16'b0000110011000110   // 51.09375
  },
  // x_re_3 = [8.171875, 3.046875, 59.5, -35.375, 31.640625, 19.5625, -26.625, 35.46875]
  {
    16'b0000001000001011,  // 8.171875
    16'b0000000011000011,  // 3.046875
    16'b0000111011100000,  // 59.5
    16'b1111011100101000,  // -35.375
    16'b0000011111101001,  // 31.640625
    16'b0000010011100100,  // 19.5625
    16'b1111100101011000,  // -26.625
    16'b0000100011011110   // 35.46875
  },
  // x_re_4 = [-16.0625, 8.8125, 38.765625, -39.78125, 53.15625, 32.9375, -50.78125, 15.078125]
  {
    16'b1111101111111100,  // -16.0625
    16'b0000001000110100,  // 8.8125
    16'b0000100110110001,  // 38.765625
    16'b1111011000001110,  // -39.78125
    16'b0000110101001010,  // 53.15625
    16'b0000100000111100,  // 32.9375
    16'b1111001101001110,  // -50.78125
    16'b0000001111000101   // 15.078125
  },
  // x_re_5 = [-52.8125, 54.46875, 31.0, -38.125, 7.8125, -27.9375, -53.34375, -10.921875]
  {
    16'b1111001011001100,  // -52.8125
    16'b0000110110011110,  // 54.46875
    16'b0000011111000000,  // 31.0
    16'b1111011001111000,  // -38.125
    16'b0000000111110100,  // 7.8125
    16'b1111100100000100,  // -27.9375
    16'b1111001010101010,  // -53.34375
    16'b1111110101000101   // -10.921875
  },
  // x_re_6 = [-39.703125, -48.28125, 49.390625, 19.171875, 2.96875, 9.0, -59.40625, 61.4375]
  {
    16'b1111011000010011,  // -39.703125
    16'b1111001111101110,  // -48.28125
    16'b0000110001011001,  // 49.390625
    16'b0000010011001011,  // 19.171875
    16'b0000000010111110,  // 2.96875
    16'b0000001001000000,  // 9.0
    16'b1111000100100110,  // -59.40625
    16'b0000111101011100   // 61.4375
  },
  // x_re_7 = [52.9375, 27.578125, -21.125, -49.078125, 43.09375, 15.875, 14.9375, 1.0]
  {
    16'b0000110100111100,  // 52.9375
    16'b0000011011100101,  // 27.578125
    16'b1111101010111000,  // -21.125
    16'b1111001110111011,  // -49.078125
    16'b0000101011000110,  // 43.09375
    16'b0000001111111000,  // 15.875
    16'b0000001110111100,  // 14.9375
    16'b0000000001000000   // 1.0
  },
  // x_re_8 = [-12.1875, 50.84375, -57.09375, -31.484375, 0.09375, -52.5625, 5.3125, 10.0625]
  {
    16'b1111110011110100,  // -12.1875
    16'b0000110010110110,  // 50.84375
    16'b1111000110111010,  // -57.09375
    16'b1111100000100001,  // -31.484375
    16'b0000000000000110,  // 0.09375
    16'b1111001011011100,  // -52.5625
    16'b0000000101010100,  // 5.3125
    16'b0000001010000100   // 10.0625
  },
  // x_re_9 = [3.734375, 1.515625, -31.609375, 55.140625, -60.796875, 19.15625, -5.578125, 11.171875]
  {
    16'b0000000011101111,  // 3.734375
    16'b0000000001100001,  // 1.515625
    16'b1111100000011001,  // -31.609375
    16'b0000110111001001,  // 55.140625
    16'b1111000011001101,  // -60.796875
    16'b0000010011001010,  // 19.15625
    16'b1111111010011011,  // -5.578125
    16'b0000001011001011   // 11.171875
  },
  // x_re_10 = [-42.578125, 24.171875, 58.359375, -6.984375, 11.421875, -21.4375, -11.5625, 30.84375]
  {
    16'b1111010101011011,  // -42.578125
    16'b0000011000001011,  // 24.171875
    16'b0000111010010111,  // 58.359375
    16'b1111111001000001,  // -6.984375
    16'b0000001011011011,  // 11.421875
    16'b1111101010100100,  // -21.4375
    16'b1111110100011100,  // -11.5625
    16'b0000011110110110   // 30.84375
  },
  // x_re_11 = [-11.046875, -61.875, -50.703125, -37.265625, -39.203125, -40.5, -30.703125, -55.484375]
  {
    16'b1111110100111101,  // -11.046875
    16'b1111000010001000,  // -61.875
    16'b1111001101010011,  // -50.703125
    16'b1111011010101111,  // -37.265625
    16'b1111011000110011,  // -39.203125
    16'b1111010111100000,  // -40.5
    16'b1111100001010011,  // -30.703125
    16'b1111001000100001   // -55.484375
  },
  // x_re_12 = [-39.0, 47.9375, -5.5, 41.75, -6.046875, -47.8125, -15.25, 40.078125]
  {
    16'b1111011001000000,  // -39.0
    16'b0000101111111100,  // 47.9375
    16'b1111111010100000,  // -5.5
    16'b0000101001110000,  // 41.75
    16'b1111111001111101,  // -6.046875
    16'b1111010000001100,  // -47.8125
    16'b1111110000110000,  // -15.25
    16'b0000101000000101   // 40.078125
  },
  // x_re_13 = [2.515625, 2.375, 29.34375, 16.78125, -36.59375, -34.0625, 37.625, -9.5625]
  {
    16'b0000000010100001,  // 2.515625
    16'b0000000010011000,  // 2.375
    16'b0000011101010110,  // 29.34375
    16'b0000010000110010,  // 16.78125
    16'b1111011011011010,  // -36.59375
    16'b1111011101111100,  // -34.0625
    16'b0000100101101000,  // 37.625
    16'b1111110110011100   // -9.5625
  },
  // x_re_14 = [-2.859375, 33.921875, 53.953125, -21.046875, 14.5625, -51.6875, -35.09375, 60.5]
  {
    16'b1111111101001001,  // -2.859375
    16'b0000100001111011,  // 33.921875
    16'b0000110101111101,  // 53.953125
    16'b1111101010111101,  // -21.046875
    16'b0000001110100100,  // 14.5625
    16'b1111001100010100,  // -51.6875
    16'b1111011100111010,  // -35.09375
    16'b0000111100100000   // 60.5
  },
  // x_re_15 = [-49.640625, 19.90625, -16.265625, -31.25, 60.171875, 20.296875, 18.390625, 45.5625]
  {
    16'b1111001110010111,  // -49.640625
    16'b0000010011111010,  // 19.90625
    16'b1111101111101111,  // -16.265625
    16'b1111100000110000,  // -31.25
    16'b0000111100001011,  // 60.171875
    16'b0000010100010011,  // 20.296875
    16'b0000010010011001,  // 18.390625
    16'b0000101101100100   // 45.5625
  },
  // x_re_16 = [55.671875, -49.640625, 59.984375, -45.78125, 38.28125, -33.546875, 27.6875, -17.59375]
  {
    16'b0000110111101011,  // 55.671875
    16'b1111001110010111,  // -49.640625
    16'b0000111011111111,  // 59.984375
    16'b1111010010001110,  // -45.78125
    16'b0000100110010010,  // 38.28125
    16'b1111011110011101,  // -33.546875
    16'b0000011011101100,  // 27.6875
    16'b1111101110011010   // -17.59375
  },
  // x_re_17 = [19.109375, -61.921875, 12.4375, -1.46875, -55.578125, 29.265625, -52.265625, -46.0]
  {
    16'b0000010011000111,  // 19.109375
    16'b1111000010000101,  // -61.921875
    16'b0000001100011100,  // 12.4375
    16'b1111111110100010,  // -1.46875
    16'b1111001000011011,  // -55.578125
    16'b0000011101010001,  // 29.265625
    16'b1111001011101111,  // -52.265625
    16'b1111010010000000   // -46.0
  },
  // x_re_18 = [-1.734375, -35.28125, -4.015625, 6.15625, 35.375, -57.671875, -44.875, 31.984375]
  {
    16'b1111111110010001,  // -1.734375
    16'b1111011100101110,  // -35.28125
    16'b1111111011111111,  // -4.015625
    16'b0000000110001010,  // 6.15625
    16'b0000100011011000,  // 35.375
    16'b1111000110010101,  // -57.671875
    16'b1111010011001000,  // -44.875
    16'b0000011111111111   // 31.984375
  },
  // x_re_19 = [38.578125, -7.21875, 59.984375, -25.9375, 51.765625, 36.609375, 50.421875, 28.296875]
  {
    16'b0000100110100101,  // 38.578125
    16'b1111111000110010,  // -7.21875
    16'b0000111011111111,  // 59.984375
    16'b1111100110000100,  // -25.9375
    16'b0000110011110001,  // 51.765625
    16'b0000100100100111,  // 36.609375
    16'b0000110010011011,  // 50.421875
    16'b0000011100010011   // 28.296875
  },
  // x_re_20 = [12.0625, 6.328125, -56.265625, 44.859375, -13.65625, 14.578125, -39.078125, 15.765625]
  {
    16'b0000001100000100,  // 12.0625
    16'b0000000110010101,  // 6.328125
    16'b1111000111101111,  // -56.265625
    16'b0000101100110111,  // 44.859375
    16'b1111110010010110,  // -13.65625
    16'b0000001110100101,  // 14.578125
    16'b1111011000111011,  // -39.078125
    16'b0000001111110001   // 15.765625
  },
  // x_re_21 = [13.515625, 52.703125, 15.078125, 57.34375, -60.03125, -23.671875, 43.234375, -48.765625]
  {
    16'b0000001101100001,  // 13.515625
    16'b0000110100101101,  // 52.703125
    16'b0000001111000101,  // 15.078125
    16'b0000111001010110,  // 57.34375
    16'b1111000011111110,  // -60.03125
    16'b1111101000010101,  // -23.671875
    16'b0000101011001111,  // 43.234375
    16'b1111001111001111   // -48.765625
  },
  // x_re_22 = [-36.875, -59.171875, 12.84375, 41.875, -53.828125, 48.203125, 35.140625, 26.234375]
  {
    16'b1111011011001000,  // -36.875
    16'b1111000100110101,  // -59.171875
    16'b0000001100110110,  // 12.84375
    16'b0000101001111000,  // 41.875
    16'b1111001010001011,  // -53.828125
    16'b0000110000001101,  // 48.203125
    16'b0000100011001001,  // 35.140625
    16'b0000011010001111   // 26.234375
  },
  // x_re_23 = [-33.765625, -62.8125, 49.34375, 46.234375, 16.984375, 6.28125, -14.359375, 34.34375]
  {
    16'b1111011110001111,  // -33.765625
    16'b1111000001001100,  // -62.8125
    16'b0000110001010110,  // 49.34375
    16'b0000101110001111,  // 46.234375
    16'b0000010000111111,  // 16.984375
    16'b0000000110010010,  // 6.28125
    16'b1111110001101001,  // -14.359375
    16'b0000100010010110   // 34.34375
  },
  // x_re_24 = [53.859375, 58.109375, 61.453125, -31.359375, -56.53125, -19.5, -63.09375, 17.140625]
  {
    16'b0000110101110111,  // 53.859375
    16'b0000111010000111,  // 58.109375
    16'b0000111101011101,  // 61.453125
    16'b1111100000101001,  // -31.359375
    16'b1111000111011110,  // -56.53125
    16'b1111101100100000,  // -19.5
    16'b1111000000111010,  // -63.09375
    16'b0000010001001001   // 17.140625
  },
  // x_re_25 = [-10.8125, -31.78125, 20.65625, 4.828125, 57.65625, 9.125, 58.734375, 55.015625]
  {
    16'b1111110101001100,  // -10.8125
    16'b1111100000001110,  // -31.78125
    16'b0000010100101010,  // 20.65625
    16'b0000000100110101,  // 4.828125
    16'b0000111001101010,  // 57.65625
    16'b0000001001001000,  // 9.125
    16'b0000111010101111,  // 58.734375
    16'b0000110111000001   // 55.015625
  },
  // x_re_26 = [44.046875, -16.515625, 39.28125, -1.21875, -47.40625, -3.4375, -2.53125, 44.65625]
  {
    16'b0000101100000011,  // 44.046875
    16'b1111101111011111,  // -16.515625
    16'b0000100111010010,  // 39.28125
    16'b1111111110110010,  // -1.21875
    16'b1111010000100110,  // -47.40625
    16'b1111111100100100,  // -3.4375
    16'b1111111101011110,  // -2.53125
    16'b0000101100101010   // 44.65625
  },
  // x_re_27 = [55.828125, 35.984375, 51.90625, -61.71875, -14.390625, -12.4375, 61.234375, -40.765625]
  {
    16'b0000110111110101,  // 55.828125
    16'b0000100011111111,  // 35.984375
    16'b0000110011111010,  // 51.90625
    16'b1111000010010010,  // -61.71875
    16'b1111110001100111,  // -14.390625
    16'b1111110011100100,  // -12.4375
    16'b0000111101001111,  // 61.234375
    16'b1111010111001111   // -40.765625
  },
  // x_re_28 = [61.546875, 30.046875, -33.0625, -27.09375, -4.859375, -35.046875, 62.296875, -41.796875]
  {
    16'b0000111101100011,  // 61.546875
    16'b0000011110000011,  // 30.046875
    16'b1111011110111100,  // -33.0625
    16'b1111100100111010,  // -27.09375
    16'b1111111011001001,  // -4.859375
    16'b1111011100111101,  // -35.046875
    16'b0000111110010011,  // 62.296875
    16'b1111010110001101   // -41.796875
  },
  // x_re_29 = [62.921875, 32.625, 36.46875, -57.515625, -20.78125, 51.75, -56.515625, 17.15625]
  {
    16'b0000111110111011,  // 62.921875
    16'b0000100000101000,  // 32.625
    16'b0000100100011110,  // 36.46875
    16'b1111000110011111,  // -57.515625
    16'b1111101011001110,  // -20.78125
    16'b0000110011110000,  // 51.75
    16'b1111000111011111,  // -56.515625
    16'b0000010001001010   // 17.15625
  },
  // x_re_30 = [10.34375, -50.953125, -6.65625, -48.546875, -34.359375, 61.75, 17.890625, -57.5625]
  {
    16'b0000001010010110,  // 10.34375
    16'b1111001101000011,  // -50.953125
    16'b1111111001010110,  // -6.65625
    16'b1111001111011101,  // -48.546875
    16'b1111011101101001,  // -34.359375
    16'b0000111101110000,  // 61.75
    16'b0000010001111001,  // 17.890625
    16'b1111000110011100   // -57.5625
  },
  // x_re_31 = [47.421875, 25.859375, 10.65625, 5.84375, 23.296875, -37.59375, 36.90625, -50.0625]
  {
    16'b0000101111011011,  // 47.421875
    16'b0000011001110111,  // 25.859375
    16'b0000001010101010,  // 10.65625
    16'b0000000101110110,  // 5.84375
    16'b0000010111010011,  // 23.296875
    16'b1111011010011010,  // -37.59375
    16'b0000100100111010,  // 36.90625
    16'b1111001101111100   // -50.0625
  },
  // x_re_32 = [-43.5, -20.25, -25.453125, -22.21875, -7.5625, -48.046875, -46.984375, 42.796875]
  {
    16'b1111010100100000,  // -43.5
    16'b1111101011110000,  // -20.25
    16'b1111100110100011,  // -25.453125
    16'b1111101001110010,  // -22.21875
    16'b1111111000011100,  // -7.5625
    16'b1111001111111101,  // -48.046875
    16'b1111010001000001,  // -46.984375
    16'b0000101010110011   // 42.796875
  },
  // x_re_33 = [-3.859375, -16.125, -53.390625, 27.015625, -51.875, 7.03125, -10.96875, -34.0625]
  {
    16'b1111111100001001,  // -3.859375
    16'b1111101111111000,  // -16.125
    16'b1111001010100111,  // -53.390625
    16'b0000011011000001,  // 27.015625
    16'b1111001100001000,  // -51.875
    16'b0000000111000010,  // 7.03125
    16'b1111110101000010,  // -10.96875
    16'b1111011101111100   // -34.0625
  },
  // x_re_34 = [22.5625, -61.546875, -14.859375, -59.15625, -5.375, 26.015625, -12.171875, 55.203125]
  {
    16'b0000010110100100,  // 22.5625
    16'b1111000010011101,  // -61.546875
    16'b1111110001001001,  // -14.859375
    16'b1111000100110110,  // -59.15625
    16'b1111111010101000,  // -5.375
    16'b0000011010000001,  // 26.015625
    16'b1111110011110101,  // -12.171875
    16'b0000110111001101   // 55.203125
  },
  // x_re_35 = [-9.59375, -50.765625, 55.28125, -43.9375, -22.0625, -63.140625, -3.328125, 23.703125]
  {
    16'b1111110110011010,  // -9.59375
    16'b1111001101001111,  // -50.765625
    16'b0000110111010010,  // 55.28125
    16'b1111010100000100,  // -43.9375
    16'b1111101001111100,  // -22.0625
    16'b1111000000110111,  // -63.140625
    16'b1111111100101011,  // -3.328125
    16'b0000010111101101   // 23.703125
  },
  // x_re_36 = [-26.96875, -19.5625, -58.625, -25.5, 3.515625, -13.90625, 37.03125, -45.453125]
  {
    16'b1111100101000010,  // -26.96875
    16'b1111101100011100,  // -19.5625
    16'b1111000101011000,  // -58.625
    16'b1111100110100000,  // -25.5
    16'b0000000011100001,  // 3.515625
    16'b1111110010000110,  // -13.90625
    16'b0000100101000010,  // 37.03125
    16'b1111010010100011   // -45.453125
  },
  // x_re_37 = [20.375, -38.78125, 31.671875, 43.765625, -33.046875, 39.453125, 56.234375, 32.5625]
  {
    16'b0000010100011000,  // 20.375
    16'b1111011001001110,  // -38.78125
    16'b0000011111101011,  // 31.671875
    16'b0000101011110001,  // 43.765625
    16'b1111011110111101,  // -33.046875
    16'b0000100111011101,  // 39.453125
    16'b0000111000001111,  // 56.234375
    16'b0000100000100100   // 32.5625
  },
  // x_re_38 = [-22.21875, 22.75, 16.578125, 21.015625, 59.734375, 52.875, 19.71875, 25.9375]
  {
    16'b1111101001110010,  // -22.21875
    16'b0000010110110000,  // 22.75
    16'b0000010000100101,  // 16.578125
    16'b0000010101000001,  // 21.015625
    16'b0000111011101111,  // 59.734375
    16'b0000110100111000,  // 52.875
    16'b0000010011101110,  // 19.71875
    16'b0000011001111100   // 25.9375
  },
  // x_re_39 = [18.84375, -28.421875, -10.203125, 46.875, -35.609375, 16.015625, -3.125, -34.578125]
  {
    16'b0000010010110110,  // 18.84375
    16'b1111100011100101,  // -28.421875
    16'b1111110101110011,  // -10.203125
    16'b0000101110111000,  // 46.875
    16'b1111011100011001,  // -35.609375
    16'b0000010000000001,  // 16.015625
    16'b1111111100111000,  // -3.125
    16'b1111011101011011   // -34.578125
  },
  // x_re_40 = [53.734375, -28.515625, 1.90625, -33.078125, 56.4375, 10.546875, -61.546875, -44.15625]
  {
    16'b0000110101101111,  // 53.734375
    16'b1111100011011111,  // -28.515625
    16'b0000000001111010,  // 1.90625
    16'b1111011110111011,  // -33.078125
    16'b0000111000011100,  // 56.4375
    16'b0000001010100011,  // 10.546875
    16'b1111000010011101,  // -61.546875
    16'b1111010011110110   // -44.15625
  },
  // x_re_41 = [55.734375, 33.890625, 29.203125, -31.3125, 30.5, 18.921875, 36.265625, 26.3125]
  {
    16'b0000110111101111,  // 55.734375
    16'b0000100001111001,  // 33.890625
    16'b0000011101001101,  // 29.203125
    16'b1111100000101100,  // -31.3125
    16'b0000011110100000,  // 30.5
    16'b0000010010111011,  // 18.921875
    16'b0000100100010001,  // 36.265625
    16'b0000011010010100   // 26.3125
  },
  // x_re_42 = [-27.03125, 46.1875, -23.796875, 19.25, 21.5, -61.703125, 63.390625, 60.890625]
  {
    16'b1111100100111110,  // -27.03125
    16'b0000101110001100,  // 46.1875
    16'b1111101000001101,  // -23.796875
    16'b0000010011010000,  // 19.25
    16'b0000010101100000,  // 21.5
    16'b1111000010010011,  // -61.703125
    16'b0000111111011001,  // 63.390625
    16'b0000111100111001   // 60.890625
  },
  // x_re_43 = [-44.265625, -6.265625, 52.734375, 39.609375, -22.15625, -35.265625, 28.234375, -56.6875]
  {
    16'b1111010011101111,  // -44.265625
    16'b1111111001101111,  // -6.265625
    16'b0000110100101111,  // 52.734375
    16'b0000100111100111,  // 39.609375
    16'b1111101001110110,  // -22.15625
    16'b1111011100101111,  // -35.265625
    16'b0000011100001111,  // 28.234375
    16'b1111000111010100   // -56.6875
  },
  // x_re_44 = [43.65625, -63.0625, -62.421875, -6.34375, 56.578125, -29.703125, -2.8125, -60.171875]
  {
    16'b0000101011101010,  // 43.65625
    16'b1111000000111100,  // -63.0625
    16'b1111000001100101,  // -62.421875
    16'b1111111001101010,  // -6.34375
    16'b0000111000100101,  // 56.578125
    16'b1111100010010011,  // -29.703125
    16'b1111111101001100,  // -2.8125
    16'b1111000011110101   // -60.171875
  },
  // x_re_45 = [-53.0, -42.234375, -27.65625, 56.53125, 20.109375, 30.46875, 1.625, -10.84375]
  {
    16'b1111001011000000,  // -53.0
    16'b1111010101110001,  // -42.234375
    16'b1111100100010110,  // -27.65625
    16'b0000111000100010,  // 56.53125
    16'b0000010100000111,  // 20.109375
    16'b0000011110011110,  // 30.46875
    16'b0000000001101000,  // 1.625
    16'b1111110101001010   // -10.84375
  },
  // x_re_46 = [60.21875, -6.609375, -5.046875, -52.0625, -29.96875, -17.9375, -53.328125, 37.09375]
  {
    16'b0000111100001110,  // 60.21875
    16'b1111111001011001,  // -6.609375
    16'b1111111010111101,  // -5.046875
    16'b1111001011111100,  // -52.0625
    16'b1111100010000010,  // -29.96875
    16'b1111101110000100,  // -17.9375
    16'b1111001010101011,  // -53.328125
    16'b0000100101000110   // 37.09375
  },
  // x_re_47 = [-52.28125, -61.234375, -35.96875, 61.84375, 1.71875, -14.828125, 3.484375, 29.265625]
  {
    16'b1111001011101110,  // -52.28125
    16'b1111000010110001,  // -61.234375
    16'b1111011100000010,  // -35.96875
    16'b0000111101110110,  // 61.84375
    16'b0000000001101110,  // 1.71875
    16'b1111110001001011,  // -14.828125
    16'b0000000011011111,  // 3.484375
    16'b0000011101010001   // 29.265625
  },
  // x_re_48 = [-8.9375, 43.0625, 59.046875, 21.546875, 61.625, -44.59375, -25.53125, 19.640625]
  {
    16'b1111110111000100,  // -8.9375
    16'b0000101011000100,  // 43.0625
    16'b0000111011000011,  // 59.046875
    16'b0000010101100011,  // 21.546875
    16'b0000111101101000,  // 61.625
    16'b1111010011011010,  // -44.59375
    16'b1111100110011110,  // -25.53125
    16'b0000010011101001   // 19.640625
  },
  // x_re_49 = [-57.796875, 61.171875, -23.140625, -17.203125, -29.515625, 38.421875, -38.984375, -13.875]
  {
    16'b1111000110001101,  // -57.796875
    16'b0000111101001011,  // 61.171875
    16'b1111101000110111,  // -23.140625
    16'b1111101110110011,  // -17.203125
    16'b1111100010011111,  // -29.515625
    16'b0000100110011011,  // 38.421875
    16'b1111011001000001,  // -38.984375
    16'b1111110010001000   // -13.875
  },
  // x_re_50 = [-20.625, -53.34375, 52.359375, 5.984375, -57.109375, -20.96875, 10.765625, -63.140625]
  {
    16'b1111101011011000,  // -20.625
    16'b1111001010101010,  // -53.34375
    16'b0000110100010111,  // 52.359375
    16'b0000000101111111,  // 5.984375
    16'b1111000110111001,  // -57.109375
    16'b1111101011000010,  // -20.96875
    16'b0000001010110001,  // 10.765625
    16'b1111000000110111   // -63.140625
  },
  // x_re_51 = [-61.796875, -30.0, 0.9375, -48.5625, -4.6875, 56.75, -17.375, 15.046875]
  {
    16'b1111000010001101,  // -61.796875
    16'b1111100010000000,  // -30.0
    16'b0000000000111100,  // 0.9375
    16'b1111001111011100,  // -48.5625
    16'b1111111011010100,  // -4.6875
    16'b0000111000110000,  // 56.75
    16'b1111101110101000,  // -17.375
    16'b0000001111000011   // 15.046875
  },
  // x_re_52 = [48.8125, 53.859375, -8.421875, 22.421875, -28.640625, 48.515625, 50.0625, -0.671875]
  {
    16'b0000110000110100,  // 48.8125
    16'b0000110101110111,  // 53.859375
    16'b1111110111100101,  // -8.421875
    16'b0000010110011011,  // 22.421875
    16'b1111100011010111,  // -28.640625
    16'b0000110000100001,  // 48.515625
    16'b0000110010000100,  // 50.0625
    16'b1111111111010101   // -0.671875
  },
  // x_re_53 = [44.5625, -2.515625, -8.359375, 33.8125, -22.59375, 46.1875, 58.265625, -44.859375]
  {
    16'b0000101100100100,  // 44.5625
    16'b1111111101011111,  // -2.515625
    16'b1111110111101001,  // -8.359375
    16'b0000100001110100,  // 33.8125
    16'b1111101001011010,  // -22.59375
    16'b0000101110001100,  // 46.1875
    16'b0000111010010001,  // 58.265625
    16'b1111010011001001   // -44.859375
  },
  // x_re_54 = [41.578125, 55.28125, 59.21875, -50.390625, 42.703125, 15.3125, -27.234375, 20.328125]
  {
    16'b0000101001100101,  // 41.578125
    16'b0000110111010010,  // 55.28125
    16'b0000111011001110,  // 59.21875
    16'b1111001101100111,  // -50.390625
    16'b0000101010101101,  // 42.703125
    16'b0000001111010100,  // 15.3125
    16'b1111100100110001,  // -27.234375
    16'b0000010100010101   // 20.328125
  },
  // x_re_55 = [22.25, 32.296875, -3.9375, -48.859375, 46.921875, 40.71875, 13.828125, -62.8125]
  {
    16'b0000010110010000,  // 22.25
    16'b0000100000010011,  // 32.296875
    16'b1111111100000100,  // -3.9375
    16'b1111001111001001,  // -48.859375
    16'b0000101110111011,  // 46.921875
    16'b0000101000101110,  // 40.71875
    16'b0000001101110101,  // 13.828125
    16'b1111000001001100   // -62.8125
  },
  // x_re_56 = [-53.59375, -21.0, 44.84375, 0.625, 52.5, 17.390625, 31.96875, -29.109375]
  {
    16'b1111001010011010,  // -53.59375
    16'b1111101011000000,  // -21.0
    16'b0000101100110110,  // 44.84375
    16'b0000000000101000,  // 0.625
    16'b0000110100100000,  // 52.5
    16'b0000010001011001,  // 17.390625
    16'b0000011111111110,  // 31.96875
    16'b1111100010111001   // -29.109375
  },
  // x_re_57 = [-20.75, -49.3125, 57.96875, 12.6875, 34.734375, -60.796875, -4.875, 45.28125]
  {
    16'b1111101011010000,  // -20.75
    16'b1111001110101100,  // -49.3125
    16'b0000111001111110,  // 57.96875
    16'b0000001100101100,  // 12.6875
    16'b0000100010101111,  // 34.734375
    16'b1111000011001101,  // -60.796875
    16'b1111111011001000,  // -4.875
    16'b0000101101010010   // 45.28125
  },
  // x_re_58 = [-50.0, 38.53125, -3.53125, -27.25, -32.59375, -11.46875, -53.140625, 19.234375]
  {
    16'b1111001110000000,  // -50.0
    16'b0000100110100010,  // 38.53125
    16'b1111111100011110,  // -3.53125
    16'b1111100100110000,  // -27.25
    16'b1111011111011010,  // -32.59375
    16'b1111110100100010,  // -11.46875
    16'b1111001010110111,  // -53.140625
    16'b0000010011001111   // 19.234375
  },
  // x_re_59 = [59.03125, -60.484375, -10.859375, -60.859375, 45.21875, 17.453125, -5.28125, -34.09375]
  {
    16'b0000111011000010,  // 59.03125
    16'b1111000011100001,  // -60.484375
    16'b1111110101001001,  // -10.859375
    16'b1111000011001001,  // -60.859375
    16'b0000101101001110,  // 45.21875
    16'b0000010001011101,  // 17.453125
    16'b1111111010101110,  // -5.28125
    16'b1111011101111010   // -34.09375
  },
  // x_re_60 = [-32.875, 19.515625, 62.609375, -17.65625, -18.609375, -41.671875, -42.734375, 23.296875]
  {
    16'b1111011111001000,  // -32.875
    16'b0000010011100001,  // 19.515625
    16'b0000111110100111,  // 62.609375
    16'b1111101110010110,  // -17.65625
    16'b1111101101011001,  // -18.609375
    16'b1111010110010101,  // -41.671875
    16'b1111010101010001,  // -42.734375
    16'b0000010111010011   // 23.296875
  },
  // x_re_61 = [28.171875, -9.8125, 58.53125, 52.25, -63.96875, -36.96875, 24.203125, 45.9375]
  {
    16'b0000011100001011,  // 28.171875
    16'b1111110110001100,  // -9.8125
    16'b0000111010100010,  // 58.53125
    16'b0000110100010000,  // 52.25
    16'b1111000000000010,  // -63.96875
    16'b1111011011000010,  // -36.96875
    16'b0000011000001101,  // 24.203125
    16'b0000101101111100   // 45.9375
  },
  // x_re_62 = [-30.75, 23.78125, 63.765625, -7.609375, 46.0, 52.546875, 46.8125, 14.828125]
  {
    16'b1111100001010000,  // -30.75
    16'b0000010111110010,  // 23.78125
    16'b0000111111110001,  // 63.765625
    16'b1111111000011001,  // -7.609375
    16'b0000101110000000,  // 46.0
    16'b0000110100100011,  // 52.546875
    16'b0000101110110100,  // 46.8125
    16'b0000001110110101   // 14.828125
  },
  // x_re_63 = [61.359375, 21.28125, 25.921875, 41.65625, 60.390625, -45.9375, -38.265625, -43.640625]
  {
    16'b0000111101010111,  // 61.359375
    16'b0000010101010010,  // 21.28125
    16'b0000011001111011,  // 25.921875
    16'b0000101001101010,  // 41.65625
    16'b0000111100011001,  // 60.390625
    16'b1111010010000100,  // -45.9375
    16'b1111011001101111,  // -38.265625
    16'b1111010100010111   // -43.640625
  }
};


logic [15 : 0] y_test_data_re [nr_of_tests_c][8] = {
  // y_re_0 = [-36.71875, -122.4375, -77.671875, 34.375, 61.0625, 34.375, -77.671875, -122.4375]
  {
    16'b1111011011010010,  // -36.71875
    16'b1110000101100100,  // -122.4375
    16'b1110110010010101,  // -77.671875
    16'b0000100010011000,  // 34.375
    16'b0000111101000100,  // 61.0625
    16'b0000100010011000,  // 34.375
    16'b1110110010010101,  // -77.671875
    16'b1110000101100100   // -122.4375
  },
  // y_re_1 = [105.6875, -20.921875, -64.078125, -128.203125, 147.84375, -128.203125, -64.078125, -20.921875]
  {
    16'b0001101001101100,  // 105.6875
    16'b1111101011000101,  // -20.921875
    16'b1110111111111011,  // -64.078125
    16'b1101111111110011,  // -128.203125
    16'b0010010011110110,  // 147.84375
    16'b1101111111110011,  // -128.203125
    16'b1110111111111011,  // -64.078125
    16'b1111101011000101   // -20.921875
  },
  // y_re_2 = [73.8125, 123.734375, 81.8125, -17.984375, -156.3125, -17.984375, 81.8125, 123.734375]
  {
    16'b0001001001110100,  // 73.8125
    16'b0001111011101111,  // 123.734375
    16'b0001010001110100,  // 81.8125
    16'b1111101110000001,  // -17.984375
    16'b1101100011101100,  // -156.3125
    16'b1111101110000001,  // -17.984375
    16'b0001010001110100,  // 81.8125
    16'b0001111011101111   // 123.734375
  },
  // y_re_3 = [95.390625, 14.71875, 6.9375, -61.65625, 49.984375, -61.65625, 6.9375, 14.71875]
  {
    16'b0001011111011001,  // 95.390625
    16'b0000001110101110,  // 14.71875
    16'b0000000110111100,  // 6.9375
    16'b1111000010010110,  // -61.65625
    16'b0000110001111111,  // 49.984375
    16'b1111000010010110,  // -61.65625
    16'b0000000110111100,  // 6.9375
    16'b0000001110101110   // 14.71875
  },
  // y_re_4 = [42.125, -47.609375, 49.109375, -90.828125, 8.03125, -90.828125, 49.109375, -47.609375]
  {
    16'b0000101010001000,  // 42.125
    16'b1111010000011001,  // -47.609375
    16'b0000110001000111,  // 49.109375
    16'b1110100101001011,  // -90.828125
    16'b0000001000000010,  // 8.03125
    16'b1110100101001011,  // -90.828125
    16'b0000110001000111,  // 49.109375
    16'b1111010000011001   // -47.609375
  },
  // y_re_5 = [-89.859375, 16.4375, -22.65625, -137.6875, -44.828125, -137.6875, -22.65625, 16.4375]
  {
    16'b1110100110001001,  // -89.859375
    16'b0000010000011100,  // 16.4375
    16'b1111101001010110,  // -22.65625
    16'b1101110110010100,  // -137.6875
    16'b1111010011001011,  // -44.828125
    16'b1101110110010100,  // -137.6875
    16'b1111101001010110,  // -22.65625
    16'b0000010000011100   // 16.4375
  },
  // y_re_6 = [-5.421875, -53.21875, -26.71875, -32.125, -88.078125, -32.125, -26.71875, -53.21875]
  {
    16'b1111111010100101,  // -5.421875
    16'b1111001010110010,  // -53.21875
    16'b1111100101010010,  // -26.71875
    16'b1111011111111000,  // -32.125
    16'b1110100111111011,  // -88.078125
    16'b1111011111111000,  // -32.125
    16'b1111100101010010,  // -26.71875
    16'b1111001010110010   // -53.21875
  },
  // y_re_7 = [85.21875, 53.28125, 102.21875, -33.59375, 94.46875, -33.59375, 102.21875, 53.28125]
  {
    16'b0001010101001110,  // 85.21875
    16'b0000110101010010,  // 53.28125
    16'b0001100110001110,  // 102.21875
    16'b1111011110011010,  // -33.59375
    16'b0001011110011110,  // 94.46875
    16'b1111011110011010,  // -33.59375
    16'b0001100110001110,  // 102.21875
    16'b0000110101010010   // 53.28125
  },
  // y_re_8 = [-87.015625, 89.625, 39.6875, -114.1875, -40.734375, -114.1875, 39.6875, 89.625]
  {
    16'b1110101000111111,  // -87.015625
    16'b0001011001101000,  // 89.625
    16'b0000100111101100,  // 39.6875
    16'b1110001101110100,  // -114.1875
    16'b1111010111010001,  // -40.734375
    16'b1110001101110100,  // -114.1875
    16'b0000100111101100,  // 39.6875
    16'b0001011001101000   // 89.625
  },
  // y_re_9 = [-7.265625, 21.21875, -19.875, 107.84375, -181.234375, 107.84375, -19.875, 21.21875]
  {
    16'b1111111000101111,  // -7.265625
    16'b0000010101001110,  // 21.21875
    16'b1111101100001000,  // -19.875
    16'b0001101011110110,  // 107.84375
    16'b1101001010110001,  // -181.234375
    16'b0001101011110110,  // 107.84375
    16'b1111101100001000,  // -19.875
    16'b0000010101001110   // 21.21875
  },
  // y_re_10 = [42.234375, 4.65625, -77.953125, -112.65625, -10.953125, -112.65625, -77.953125, 4.65625]
  {
    16'b0000101010001111,  // 42.234375
    16'b0000000100101010,  // 4.65625
    16'b1110110010000011,  // -77.953125
    16'b1110001111010110,  // -112.65625
    16'b1111110101000011,  // -10.953125
    16'b1110001111010110,  // -112.65625
    16'b1110110010000011,  // -77.953125
    16'b0000000100101010   // 4.65625
  },
  // y_re_11 = [-326.78125, 0.328125, 31.15625, 55.984375, 63.46875, 55.984375, 31.15625, 0.328125]
  {
    16'b1010111001001110,  // -326.78125
    16'b0000000000010101,  // 0.328125
    16'b0000011111001010,  // 31.15625
    16'b0000110111111111,  // 55.984375
    16'b0000111111011110,  // 63.46875
    16'b0000110111111111,  // 55.984375
    16'b0000011111001010,  // 31.15625
    16'b0000000000010101   // 0.328125
  },
  // y_re_12 = [16.15625, 33.1875, -24.296875, -99.09375, -147.75, -99.09375, -24.296875, 33.1875]
  {
    16'b0000010000001010,  // 16.15625
    16'b0000100001001100,  // 33.1875
    16'b1111100111101101,  // -24.296875
    16'b1110011100111010,  // -99.09375
    16'b1101101100010000,  // -147.75
    16'b1110011100111010,  // -99.09375
    16'b1111100111101101,  // -24.296875
    16'b0000100001001100   // 33.1875
  },
  // y_re_13 = [8.421875, 46.203125, -101.046875, 32.015625, 57.359375, 32.015625, -101.046875, 46.203125]
  {
    16'b0000001000011011,  // 8.421875
    16'b0000101110001101,  // 46.203125
    16'b1110011010111101,  // -101.046875
    16'b0000100000000001,  // 32.015625
    16'b0000111001010111,  // 57.359375
    16'b0000100000000001,  // 32.015625
    16'b1110011010111101,  // -101.046875
    16'b0000101110001101   // 46.203125
  },
  // y_re_14 = [52.25, 100.109375, -7.15625, -134.953125, 8.875, -134.953125, -7.15625, 100.109375]
  {
    16'b0000110100010000,  // 52.25
    16'b0001100100000111,  // 100.109375
    16'b1111111000110110,  // -7.15625
    16'b1101111001000011,  // -134.953125
    16'b0000001000111000,  // 8.875
    16'b1101111001000011,  // -134.953125
    16'b1111111000110110,  // -7.15625
    16'b0001100100000111   // 100.109375
  },
  // y_re_15 = [67.171875, -56.09375, 8.40625, -163.53125, -41.859375, -163.53125, 8.40625, -56.09375]
  {
    16'b0001000011001011,  // 67.171875
    16'b1111000111111010,  // -56.09375
    16'b0000001000011010,  // 8.40625
    16'b1101011100011110,  // -163.53125
    16'b1111010110001001,  // -41.859375
    16'b1101011100011110,  // -163.53125
    16'b0000001000011010,  // 8.40625
    16'b1111000111111010   // -56.09375
  },
  // y_re_16 = [35.0625, 25.890625, 6.28125, 8.890625, 328.1875, 8.890625, 6.28125, 25.890625]
  {
    16'b0000100011000100,  // 35.0625
    16'b0000011001111001,  // 25.890625
    16'b0000000110010010,  // 6.28125
    16'b0000001000111001,  // 8.890625
    16'b0101001000001100,  // 328.1875
    16'b0000001000111001,  // 8.890625
    16'b0000000110010010,  // 6.28125
    16'b0000011001111001   // 25.890625
  },
  // y_re_17 = [-156.421875, -20.734375, 3.359375, 170.109375, 3.828125, 170.109375, 3.359375, -20.734375]
  {
    16'b1101100011100101,  // -156.421875
    16'b1111101011010001,  // -20.734375
    16'b0000000011010111,  // 3.359375
    16'b0010101010000111,  // 170.109375
    16'b0000000011110101,  // 3.828125
    16'b0010101010000111,  // 170.109375
    16'b0000000011010111,  // 3.359375
    16'b1111101011010001   // -20.734375
  },
  // y_re_18 = [-70.0625, -3.21875, 82.53125, -71.0, 39.5625, -71.0, 82.53125, -3.21875]
  {
    16'b1110111001111100,  // -70.0625
    16'b1111111100110010,  // -3.21875
    16'b0001010010100010,  // 82.53125
    16'b1110111001000000,  // -71.0
    16'b0000100111100100,  // 39.5625
    16'b1110111001000000,  // -71.0
    16'b0001010010100010,  // 82.53125
    16'b1111111100110010   // -3.21875
  },
  // y_re_19 = [232.5, -5.875, -20.0625, -20.5, 169.0, -20.5, -20.0625, -5.875]
  {
    16'b0011101000100000,  // 232.5
    16'b1111111010001000,  // -5.875
    16'b1111101011111100,  // -20.0625
    16'b1111101011100000,  // -20.5
    16'b0010101001000000,  // 169.0
    16'b1111101011100000,  // -20.5
    16'b1111101011111100,  // -20.0625
    16'b1111111010001000   // -5.875
  },
  // y_re_20 = [-15.40625, -0.53125, 93.75, 51.96875, -178.46875, 51.96875, 93.75, -0.53125]
  {
    16'b1111110000100110,  // -15.40625
    16'b1111111111011110,  // -0.53125
    16'b0001011101110000,  // 93.75
    16'b0000110011111110,  // 51.96875
    16'b1101001101100010,  // -178.46875
    16'b0000110011111110,  // 51.96875
    16'b0001011101110000,  // 93.75
    16'b1111111111011110   // -0.53125
  },
  // y_re_21 = [49.40625, 52.640625, -104.828125, 94.453125, -25.8125, 94.453125, -104.828125, 52.640625]
  {
    16'b0000110001011010,  // 49.40625
    16'b0000110100101001,  // 52.640625
    16'b1110010111001011,  // -104.828125
    16'b0001011110011101,  // 94.453125
    16'b1111100110001100,  // -25.8125
    16'b0001011110011101,  // 94.453125
    16'b1110010111001011,  // -104.828125
    16'b0000110100101001   // 52.640625
  },
  // y_re_22 = [14.421875, -69.53125, -138.6875, 103.4375, -99.859375, 103.4375, -138.6875, -69.53125]
  {
    16'b0000001110011011,  // 14.421875
    16'b1110111010011110,  // -69.53125
    16'b1101110101010100,  // -138.6875
    16'b0001100111011100,  // 103.4375
    16'b1110011100001001,  // -99.859375
    16'b0001100111011100,  // 103.4375
    16'b1101110101010100,  // -138.6875
    16'b1110111010011110   // -69.53125
  },
  // y_re_23 = [42.25, -107.6875, -51.765625, 6.1875, -5.84375, 6.1875, -51.765625, -107.6875]
  {
    16'b0000101010010000,  // 42.25
    16'b1110010100010100,  // -107.6875
    16'b1111001100001111,  // -51.765625
    16'b0000000110001100,  // 6.1875
    16'b1111111010001010,  // -5.84375
    16'b0000000110001100,  // 6.1875
    16'b1111001100001111,  // -51.765625
    16'b1110010100010100   // -107.6875
  },
  // y_re_24 = [20.078125, 199.046875, -1.03125, 21.734375, -28.703125, 21.734375, -1.03125, 199.046875]
  {
    16'b0000010100000101,  // 20.078125
    16'b0011000111000011,  // 199.046875
    16'b1111111110111110,  // -1.03125
    16'b0000010101101111,  // 21.734375
    16'b1111100011010011,  // -28.703125
    16'b0000010101101111,  // 21.734375
    16'b1111111110111110,  // -1.03125
    16'b0011000111000011   // 199.046875
  },
  // y_re_25 = [163.421875, -61.953125, -32.546875, -74.984375, 89.046875, -74.984375, -32.546875, -61.953125]
  {
    16'b0010100011011011,  // 163.421875
    16'b1111000010000011,  // -61.953125
    16'b1111011111011101,  // -32.546875
    16'b1110110101000001,  // -74.984375
    16'b0001011001000011,  // 89.046875
    16'b1110110101000001,  // -74.984375
    16'b1111011111011101,  // -32.546875
    16'b1111000010000011   // -61.953125
  },
  // y_re_26 = [56.875, 114.5, -40.109375, 68.40625, 9.90625, 68.40625, -40.109375, 114.5]
  {
    16'b0000111000111000,  // 56.875
    16'b0001110010100000,  // 114.5
    16'b1111010111111001,  // -40.109375
    16'b0001000100011010,  // 68.40625
    16'b0000001001111010,  // 9.90625
    16'b0001000100011010,  // 68.40625
    16'b1111010111111001,  // -40.109375
    16'b0001110010100000   // 114.5
  },
  // y_re_27 = [75.640625, 118.984375, -71.703125, 21.453125, 233.515625, 21.453125, -71.703125, 118.984375]
  {
    16'b0001001011101001,  // 75.640625
    16'b0001110110111111,  // 118.984375
    16'b1110111000010011,  // -71.703125
    16'b0000010101011101,  // 21.453125
    16'b0011101001100001,  // 233.515625
    16'b0000010101011101,  // 21.453125
    16'b1110111000010011,  // -71.703125
    16'b0001110110111111   // 118.984375
  },
  // y_re_28 = [12.03125, 101.828125, 27.453125, 30.984375, 159.8125, 30.984375, 27.453125, 101.828125]
  {
    16'b0000001100000010,  // 12.03125
    16'b0001100101110101,  // 101.828125
    16'b0000011011011101,  // 27.453125
    16'b0000011110111111,  // 30.984375
    16'b0010011111110100,  // 159.8125
    16'b0000011110111111,  // 30.984375
    16'b0000011011011101,  // 27.453125
    16'b0001100101110101   // 101.828125
  },
  // y_re_29 = [66.109375, 122.75, 62.1875, 44.65625, -21.921875, 44.65625, 62.1875, 122.75]
  {
    16'b0001000010000111,  // 66.109375
    16'b0001111010110000,  // 122.75
    16'b0000111110001100,  // 62.1875
    16'b0000101100101010,  // 44.65625
    16'b1111101010000101,  // -21.921875
    16'b0000101100101010,  // 44.65625
    16'b0000111110001100,  // 62.1875
    16'b0001111010110000   // 122.75
  },
  // y_re_30 = [-108.09375, -40.875, -35.25, 130.28125, 82.53125, 130.28125, -35.25, -40.875]
  {
    16'b1110010011111010,  // -108.09375
    16'b1111010111001000,  // -40.875
    16'b1111011100110000,  // -35.25
    16'b0010000010010010,  // 130.28125
    16'b0001010010100010,  // 82.53125
    16'b0010000010010010,  // 130.28125
    16'b1111011100110000,  // -35.25
    16'b1111010111001000   // -40.875
  },
  // y_re_31 = [62.328125, 29.421875, 23.15625, 18.828125, 174.234375, 18.828125, 23.15625, 29.421875]
  {
    16'b0000111110010101,  // 62.328125
    16'b0000011101011011,  // 29.421875
    16'b0000010111001010,  // 23.15625
    16'b0000010010110101,  // 18.828125
    16'b0010101110001111,  // 174.234375
    16'b0000010010110101,  // 18.828125
    16'b0000010111001010,  // 23.15625
    16'b0000011101011011   // 29.421875
  },
  // y_re_32 = [-171.21875, 29.3125, 21.375, -101.1875, -75.78125, -101.1875, 21.375, 29.3125]
  {
    16'b1101010100110010,  // -171.21875
    16'b0000011101010100,  // 29.3125
    16'b0000010101011000,  // 21.375
    16'b1110011010110100,  // -101.1875
    16'b1110110100001110,  // -75.78125
    16'b1110011010110100,  // -101.1875
    16'b0000010101011000,  // 21.375
    16'b0000011101010100   // 29.3125
  },
  // y_re_33 = [-136.234375, -11.203125, 8.625, 107.234375, -103.953125, 107.234375, 8.625, -11.203125]
  {
    16'b1101110111110001,  // -136.234375
    16'b1111110100110011,  // -11.203125
    16'b0000001000101000,  // 8.625
    16'b0001101011001111,  // 107.234375
    16'b1110011000000011,  // -103.953125
    16'b0001101011001111,  // 107.234375
    16'b0000001000101000,  // 8.625
    16'b1111110100110011   // -11.203125
  },
  // y_re_34 = [-49.328125, 46.765625, 44.21875, 9.109375, 29.640625, 9.109375, 44.21875, 46.765625]
  {
    16'b1111001110101011,  // -49.328125
    16'b0000101110110001,  // 46.765625
    16'b0000101100001110,  // 44.21875
    16'b0000001001000111,  // 9.109375
    16'b0000011101101001,  // 29.640625
    16'b0000001001000111,  // 9.109375
    16'b0000101100001110,  // 44.21875
    16'b0000101110110001   // 46.765625
  },
  // y_re_35 = [-113.84375, 68.71875, -83.609375, -43.78125, 154.4375, -43.78125, -83.609375, 68.71875]
  {
    16'b1110001110001010,  // -113.84375
    16'b0001000100101110,  // 68.71875
    16'b1110101100011001,  // -83.609375
    16'b1111010100001110,  // -43.78125
    16'b0010011010011100,  // 154.4375
    16'b1111010100001110,  // -43.78125
    16'b1110101100011001,  // -83.609375
    16'b0001000100101110   // 68.71875
  },
  // y_re_36 = [-149.46875, -48.484375, -1.859375, -12.484375, 59.375, -12.484375, -1.859375, -48.484375]
  {
    16'b1101101010100010,  // -149.46875
    16'b1111001111100001,  // -48.484375
    16'b1111111110001001,  // -1.859375
    16'b1111110011100001,  // -12.484375
    16'b0000111011011000,  // 59.375
    16'b1111110011100001,  // -12.484375
    16'b1111111110001001,  // -1.859375
    16'b1111001111100001   // -48.484375
  },
  // y_re_37 = [152.234375, -9.453125, -100.578125, 116.296875, -1.765625, 116.296875, -100.578125, -9.453125]
  {
    16'b0010011000001111,  // 152.234375
    16'b1111110110100011,  // -9.453125
    16'b1110011011011011,  // -100.578125
    16'b0001110100010011,  // 116.296875
    16'b1111111110001111,  // -1.765625
    16'b0001110100010011,  // 116.296875
    16'b1110011011011011,  // -100.578125
    16'b1111110110100011   // -9.453125
  },
  // y_re_38 = [196.390625, -99.671875, 1.21875, -64.234375, -48.765625, -64.234375, 1.21875, -99.671875]
  {
    16'b0011000100011001,  // 196.390625
    16'b1110011100010101,  // -99.671875
    16'b0000000001001110,  // 1.21875
    16'b1110111111110001,  // -64.234375
    16'b1111001111001111,  // -48.765625
    16'b1110111111110001,  // -64.234375
    16'b0000000001001110,  // 1.21875
    16'b1110011100010101   // -99.671875
  },
  // y_re_39 = [-30.203125, -34.0625, -3.4375, 142.96875, -29.984375, 142.96875, -3.4375, -34.0625]
  {
    16'b1111100001110011,  // -30.203125
    16'b1111011101111100,  // -34.0625
    16'b1111111100100100,  // -3.4375
    16'b0010001110111110,  // 142.96875
    16'b1111100010000001,  // -29.984375
    16'b0010001110111110,  // 142.96875
    16'b1111111100100100,  // -3.4375
    16'b1111011101111100   // -34.0625
  },
  // y_re_40 = [-44.671875, -37.953125, 169.8125, 32.546875, 145.734375, 32.546875, 169.8125, -37.953125]
  {
    16'b1111010011010101,  // -44.671875
    16'b1111011010000011,  // -37.953125
    16'b0010101001110100,  // 169.8125
    16'b0000100000100011,  // 32.546875
    16'b0010010001101111,  // 145.734375
    16'b0000100000100011,  // 32.546875
    16'b0010101001110100,  // 169.8125
    16'b1111011010000011   // -37.953125
  },
  // y_re_41 = [199.515625, 76.265625, 20.765625, -25.796875, 103.890625, -25.796875, 20.765625, 76.265625]
  {
    16'b0011000111100001,  // 199.515625
    16'b0001001100010001,  // 76.265625
    16'b0000010100110001,  // 20.765625
    16'b1111100110001101,  // -25.796875
    16'b0001100111111001,  // 103.890625
    16'b1111100110001101,  // -25.796875
    16'b0000010100110001,  // 20.765625
    16'b0001001100010001   // 76.265625
  },
  // y_re_42 = [98.6875, 56.59375, -45.125, -153.65625, -30.5625, -153.65625, -45.125, 56.59375]
  {
    16'b0001100010101100,  // 98.6875
    16'b0000111000100110,  // 56.59375
    16'b1111010010111000,  // -45.125
    16'b1101100110010110,  // -153.65625
    16'b1111100001011100,  // -30.5625
    16'b1101100110010110,  // -153.65625
    16'b1111010010111000,  // -45.125
    16'b0000111000100110   // 56.59375
  },
  // y_re_43 = [-44.0625, -69.421875, -147.390625, 25.203125, 73.15625, 25.203125, -147.390625, -69.421875]
  {
    16'b1111010011111100,  // -44.0625
    16'b1110111010100101,  // -69.421875
    16'b1101101100100111,  // -147.390625
    16'b0000011001001101,  // 25.203125
    16'b0001001001001010,  // 73.15625
    16'b0000011001001101,  // 25.203125
    16'b1101101100100111,  // -147.390625
    16'b1110111010100101   // -69.421875
  },
  // y_re_44 = [-124.28125, -74.21875, 165.46875, 48.375, 194.28125, 48.375, 165.46875, -74.21875]
  {
    16'b1110000011101110,  // -124.28125
    16'b1110110101110010,  // -74.21875
    16'b0010100101011110,  // 165.46875
    16'b0000110000011000,  // 48.375
    16'b0011000010010010,  // 194.28125
    16'b0000110000011000,  // 48.375
    16'b0010100101011110,  // 165.46875
    16'b1110110101110010   // -74.21875
  },
  // y_re_45 = [-25.0, -171.59375, -6.859375, 25.375, -92.84375, 25.375, -6.859375, -171.59375]
  {
    16'b1111100111000000,  // -25.0
    16'b1101010100011010,  // -171.59375
    16'b1111111001001001,  // -6.859375
    16'b0000011001011000,  // 25.375
    16'b1110100011001010,  // -92.84375
    16'b0000011001011000,  // 25.375
    16'b1111111001001001,  // -6.859375
    16'b1101010100011010   // -171.59375
  },
  // y_re_46 = [-67.640625, 160.828125, 88.625, 19.546875, 11.390625, 19.546875, 88.625, 160.828125]
  {
    16'b1110111100010111,  // -67.640625
    16'b0010100000110101,  // 160.828125
    16'b0001011000101000,  // 88.625
    16'b0000010011100011,  // 19.546875
    16'b0000001011011001,  // 11.390625
    16'b0000010011100011,  // 19.546875
    16'b0001011000101000,  // 88.625
    16'b0010100000110101   // 160.828125
  },
  // y_re_47 = [-68.0, -109.53125, -18.078125, 1.53125, -98.09375, 1.53125, -18.078125, -109.53125]
  {
    16'b1110111100000000,  // -68.0
    16'b1110010010011110,  // -109.53125
    16'b1111101101111011,  // -18.078125
    16'b0000000001100010,  // 1.53125
    16'b1110011101111010,  // -98.09375
    16'b0000000001100010,  // 1.53125
    16'b1111101101111011,  // -18.078125
    16'b1110010010011110   // -109.53125
  },
  // y_re_48 = [125.859375, -10.28125, 19.171875, -130.84375, 46.546875, -130.84375, 19.171875, -10.28125]
  {
    16'b0001111101110111,  // 125.859375
    16'b1111110101101110,  // -10.28125
    16'b0000010011001011,  // 19.171875
    16'b1101111101001010,  // -130.84375
    16'b0000101110100011,  // 46.546875
    16'b1101111101001010,  // -130.84375
    16'b0000010011001011,  // 19.171875
    16'b1111110101101110   // -10.28125
  },
  // y_re_49 = [-80.921875, -9.953125, -25.1875, -46.609375, -217.953125, -46.609375, -25.1875, -9.953125]
  {
    16'b1110101111000101,  // -80.921875
    16'b1111110110000011,  // -9.953125
    16'b1111100110110100,  // -25.1875
    16'b1111010001011001,  // -46.609375
    16'b1100100110000011,  // -217.953125
    16'b1111010001011001,  // -46.609375
    16'b1111100110110100,  // -25.1875
    16'b1111110110000011   // -9.953125
  },
  // y_re_50 = [-146.078125, -34.875, -140.859375, 107.84375, 116.859375, 107.84375, -140.859375, -34.875]
  {
    16'b1101101101111011,  // -146.078125
    16'b1111011101001000,  // -34.875
    16'b1101110011001001,  // -140.859375
    16'b0001101011110110,  // 107.84375
    16'b0001110100110111,  // 116.859375
    16'b0001101011110110,  // 107.84375
    16'b1101110011001001,  // -140.859375
    16'b1111011101001000   // -34.875
  },
  // y_re_51 = [-89.6875, -73.375, -50.046875, -40.84375, -76.15625, -40.84375, -50.046875, -73.375]
  {
    16'b1110100110010100,  // -89.6875
    16'b1110110110101000,  // -73.375
    16'b1111001101111101,  // -50.046875
    16'b1111010111001010,  // -40.84375
    16'b1110110011110110,  // -76.15625
    16'b1111010111001010,  // -40.84375
    16'b1111001101111101,  // -50.046875
    16'b1110110110101000   // -73.375
  },
  // y_re_52 = [185.9375, 64.984375, -21.46875, 89.921875, -62.3125, 89.921875, -21.46875, 64.984375]
  {
    16'b0010111001111100,  // 185.9375
    16'b0001000000111111,  // 64.984375
    16'b1111101010100010,  // -21.46875
    16'b0001011001111011,  // 89.921875
    16'b1111000001101100,  // -62.3125
    16'b0001011001111011,  // 89.921875
    16'b1111101010100010,  // -21.46875
    16'b0001000000111111   // 64.984375
  },
  // y_re_53 = [104.5, -22.390625, -27.9375, 156.703125, 39.25, 156.703125, -27.9375, -22.390625]
  {
    16'b0001101000100000,  // 104.5
    16'b1111101001100111,  // -22.390625
    16'b1111100100000100,  // -27.9375
    16'b0010011100101101,  // 156.703125
    16'b0000100111010000,  // 39.25
    16'b0010011100101101,  // 156.703125
    16'b1111100100000100,  // -27.9375
    16'b1111101001100111   // -22.390625
  },
  // y_re_54 = [156.796875, 76.6875, 52.296875, -78.9375, 75.734375, -78.9375, 52.296875, 76.6875]
  {
    16'b0010011100110011,  // 156.796875
    16'b0001001100101100,  // 76.6875
    16'b0000110100010011,  // 52.296875
    16'b1110110001000100,  // -78.9375
    16'b0001001011101111,  // 75.734375
    16'b1110110001000100,  // -78.9375
    16'b0000110100010011,  // 52.296875
    16'b0001001100101100   // 76.6875
  },
  // y_re_55 = [40.40625, -40.390625, 59.28125, -8.953125, 117.71875, -8.953125, 59.28125, -40.390625]
  {
    16'b0000101000011010,  // 40.40625
    16'b1111010111100111,  // -40.390625
    16'b0000111011010010,  // 59.28125
    16'b1111110111000011,  // -8.953125
    16'b0001110101101110,  // 117.71875
    16'b1111110111000011,  // -8.953125
    16'b0000111011010010,  // 59.28125
    16'b1111010111100111   // -40.390625
  },
  // y_re_56 = [43.625, -153.984375, -77.90625, -58.203125, 107.8125, -58.203125, -77.90625, -153.984375]
  {
    16'b0000101011101000,  // 43.625
    16'b1101100110000001,  // -153.984375
    16'b1110110010000110,  // -77.90625
    16'b1111000101110011,  // -58.203125
    16'b0001101011110100,  // 107.8125
    16'b1111000101110011,  // -58.203125
    16'b1110110010000110,  // -77.90625
    16'b1101100110000001   // -153.984375
  },
  // y_re_57 = [14.9375, -24.5, -39.109375, -86.46875, 119.21875, -86.46875, -39.109375, -24.5]
  {
    16'b0000001110111100,  // 14.9375
    16'b1111100111100000,  // -24.5
    16'b1111011000111001,  // -39.109375
    16'b1110101001100010,  // -86.46875
    16'b0001110111001110,  // 119.21875
    16'b1110101001100010,  // -86.46875
    16'b1111011000111001,  // -39.109375
    16'b1111100111100000   // -24.5
  },
  // y_re_58 = [-120.21875, 50.421875, -25.921875, -85.234375, -158.3125, -85.234375, -25.921875, 50.421875]
  {
    16'b1110000111110010,  // -120.21875
    16'b0000110010011011,  // 50.421875
    16'b1111100110000101,  // -25.921875
    16'b1110101010110001,  // -85.234375
    16'b1101100001101100,  // -158.3125
    16'b1110101010110001,  // -85.234375
    16'b1111100110000101,  // -25.921875
    16'b0000110010011011   // 50.421875
  },
  // y_re_59 = [-49.875, -22.15625, 120.390625, 49.78125, 226.09375, 49.78125, 120.390625, -22.15625]
  {
    16'b1111001110001000,  // -49.875
    16'b1111101001110110,  // -22.15625
    16'b0001111000011001,  // 120.390625
    16'b0000110001110010,  // 49.78125
    16'b0011100010000110,  // 226.09375
    16'b0000110001110010,  // 49.78125
    16'b0001111000011001,  // 120.390625
    16'b1111101001110110   // -22.15625
  },
  // y_re_60 = [-48.125, 57.546875, -71.359375, -86.078125, -15.09375, -86.078125, -71.359375, 57.546875]
  {
    16'b1111001111111000,  // -48.125
    16'b0000111001100011,  // 57.546875
    16'b1110111000101001,  // -71.359375
    16'b1110101001111011,  // -86.078125
    16'b1111110000111010,  // -15.09375
    16'b1110101001111011,  // -86.078125
    16'b1110111000101001,  // -71.359375
    16'b0000111001100011   // 57.546875
  },
  // y_re_61 = [98.34375, 106.78125, -118.53125, 77.5, -4.46875, 77.5, -118.53125, 106.78125]
  {
    16'b0001100010010110,  // 98.34375
    16'b0001101010110010,  // 106.78125
    16'b1110001001011110,  // -118.53125
    16'b0001001101100000,  // 77.5
    16'b1111111011100010,  // -4.46875
    16'b0001001101100000,  // 77.5
    16'b1110001001011110,  // -118.53125
    16'b0001101010110010   // 106.78125
  },
  // y_re_62 = [209.375, -81.1875, -95.328125, -72.3125, 42.28125, -72.3125, -95.328125, -81.1875]
  {
    16'b0011010001011000,  // 209.375
    16'b1110101110110100,  // -81.1875
    16'b1110100000101011,  // -95.328125
    16'b1110110111101100,  // -72.3125
    16'b0000101010010010,  // 42.28125
    16'b1110110111101100,  // -72.3125
    16'b1110100000101011,  // -95.328125
    16'b1110101110110100   // -81.1875
  },
  // y_re_63 = [82.765625, -11.734375, 134.09375, 13.671875, 136.046875, 13.671875, 134.09375, -11.734375]
  {
    16'b0001010010110001,  // 82.765625
    16'b1111110100010001,  // -11.734375
    16'b0010000110000110,  // 134.09375
    16'b0000001101101011,  // 13.671875
    16'b0010001000000011,  // 136.046875
    16'b0000001101101011,  // 13.671875
    16'b0010000110000110,  // 134.09375
    16'b1111110100010001   // -11.734375
  }
};


logic [15 : 0] y_test_data_im [nr_of_tests_c][8] = {
  // y_im_0 = [0.0, -34.59375, 34.078125, -35.25, 0.0, 35.25, -34.078125, 34.59375]
  {
    16'b0000000000000000,  // 0.0
    16'b1111011101011010,  // -34.59375
    16'b0000100010000101,  // 34.078125
    16'b1111011100110000,  // -35.25
    16'b0000000000000000,  // 0.0
    16'b0000100011010000,  // 35.25
    16'b1111011101111011,  // -34.078125
    16'b0000100010100110   // 34.59375
  },
  // y_im_1 = [0.0, -15.96875, -8.765625, -65.0, 0.0, 65.0, 8.765625, 15.96875]
  {
    16'b0000000000000000,  // 0.0
    16'b1111110000000010,  // -15.96875
    16'b1111110111001111,  // -8.765625
    16'b1110111111000000,  // -65.0
    16'b0000000000000000,  // 0.0
    16'b0001000001000000,  // 65.0
    16'b0000001000110001,  // 8.765625
    16'b0000001111111110   // 15.96875
  },
  // y_im_2 = [0.0, 103.5, -95.78125, 15.0625, 0.0, -15.0625, 95.78125, -103.5]
  {
    16'b0000000000000000,  // 0.0
    16'b0001100111100000,  // 103.5
    16'b1110100000001110,  // -95.78125
    16'b0000001111000100,  // 15.0625
    16'b0000000000000000,  // 0.0
    16'b1111110000111100,  // -15.0625
    16'b0001011111110010,  // 95.78125
    16'b1110011000100000   // -103.5
  },
  // y_im_3 = [0.0, -24.703125, -22.515625, 147.546875, 0.0, -147.546875, 22.515625, 24.703125]
  {
    16'b0000000000000000,  // 0.0
    16'b1111100111010011,  // -24.703125
    16'b1111101001011111,  // -22.515625
    16'b0010010011100011,  // 147.546875
    16'b0000000000000000,  // 0.0
    16'b1101101100011101,  // -147.546875
    16'b0000010110100001,  // 22.515625
    16'b0000011000101101   // 24.703125
  },
  // y_im_4 = [0.0, -34.015625, -66.453125, 145.078125, 0.0, -145.078125, 66.453125, 34.015625]
  {
    16'b0000000000000000,  // 0.0
    16'b1111011101111111,  // -34.015625
    16'b1110111101100011,  // -66.453125
    16'b0010010001000101,  // 145.078125
    16'b0000000000000000,  // 0.0
    16'b1101101110111011,  // -145.078125
    16'b0001000010011101,  // 66.453125
    16'b0000100010000001   // 34.015625
  },
  // y_im_5 = [0.0, -123.15625, -75.578125, 45.53125, 0.0, -45.53125, 75.578125, 123.15625]
  {
    16'b0000000000000000,  // 0.0
    16'b1110000100110110,  // -123.15625
    16'b1110110100011011,  // -75.578125
    16'b0000101101100010,  // 45.53125
    16'b0000000000000000,  // 0.0
    16'b1111010010011110,  // -45.53125
    16'b0001001011100101,  // 75.578125
    16'b0001111011001010   // 123.15625
  },
  // y_im_6 = [0.0, -38.8125, 119.890625, 178.78125, 0.0, -178.78125, -119.890625, 38.8125]
  {
    16'b0000000000000000,  // 0.0
    16'b1111011001001100,  // -38.8125
    16'b0001110111111001,  // 119.890625
    16'b0010110010110010,  // 178.78125
    16'b0000000000000000,  // 0.0
    16'b1101001101001110,  // -178.78125
    16'b1110001000000111,  // -119.890625
    16'b0000100110110100   // 38.8125
  },
  // y_im_7 = [0.0, 63.03125, -91.53125, -9.09375, 0.0, 9.09375, 91.53125, -63.03125]
  {
    16'b0000000000000000,  // 0.0
    16'b0000111111000010,  // 63.03125
    16'b1110100100011110,  // -91.53125
    16'b1111110110111010,  // -9.09375
    16'b0000000000000000,  // 0.0
    16'b0000001001000110,  // 9.09375
    16'b0001011011100010,  // 91.53125
    16'b1111000000111110   // -63.03125
  },
  // y_im_8 = [0.0, 18.921875, -19.703125, -105.890625, 0.0, 105.890625, 19.703125, -18.921875]
  {
    16'b0000000000000000,  // 0.0
    16'b0000010010111011,  // 18.921875
    16'b1111101100010011,  // -19.703125
    16'b1110010110000111,  // -105.890625
    16'b0000000000000000,  // 0.0
    16'b0001101001111001,  // 105.890625
    16'b0000010011101101,  // 19.703125
    16'b1111101101000101   // -18.921875
  },
  // y_im_9 = [0.0, 7.53125, 45.640625, -44.53125, 0.0, 44.53125, -45.640625, -7.53125]
  {
    16'b0000000000000000,  // 0.0
    16'b0000000111100010,  // 7.53125
    16'b0000101101101001,  // 45.640625
    16'b1111010011011110,  // -44.53125
    16'b0000000000000000,  // 0.0
    16'b0000101100100010,  // 44.53125
    16'b1111010010010111,  // -45.640625
    16'b1111111000011110   // -7.53125
  },
  // y_im_10 = [0.0, -75.390625, 21.125, 64.453125, 0.0, -64.453125, -21.125, 75.390625]
  {
    16'b0000000000000000,  // 0.0
    16'b1110110100100111,  // -75.390625
    16'b0000010101001000,  // 21.125
    16'b0001000000011101,  // 64.453125
    16'b0000000000000000,  // 0.0
    16'b1110111111100011,  // -64.453125
    16'b1111101010111000,  // -21.125
    16'b0001001011011001   // 75.390625
  },
  // y_im_11 = [0.0, 22.21875, 9.625, -17.78125, 0.0, 17.78125, -9.625, -22.21875]
  {
    16'b0000000000000000,  // 0.0
    16'b0000010110001110,  // 22.21875
    16'b0000001001101000,  // 9.625
    16'b1111101110001110,  // -17.78125
    16'b0000000000000000,  // 0.0
    16'b0000010001110010,  // 17.78125
    16'b1111110110011000,  // -9.625
    16'b1111101001110010   // -22.21875
  },
  // y_im_12 = [0.0, -78.234375, 81.703125, -58.734375, 0.0, 58.734375, -81.703125, 78.234375]
  {
    16'b0000000000000000,  // 0.0
    16'b1110110001110001,  // -78.234375
    16'b0001010001101101,  // 81.703125
    16'b1111000101010001,  // -58.734375
    16'b0000000000000000,  // 0.0
    16'b0000111010101111,  // 58.734375
    16'b1110101110010011,  // -81.703125
    16'b0001001110001111   // 78.234375
  },
  // y_im_13 = [0.0, -35.859375, 38.90625, -52.421875, 0.0, 52.421875, -38.90625, 35.859375]
  {
    16'b0000000000000000,  // 0.0
    16'b1111011100001001,  // -35.859375
    16'b0000100110111010,  // 38.90625
    16'b1111001011100101,  // -52.421875
    16'b0000000000000000,  // 0.0
    16'b0000110100011011,  // 52.421875
    16'b1111011001000110,  // -38.90625
    16'b0000100011110111   // 35.859375
  },
  // y_im_14 = [0.0, -91.890625, 57.21875, 86.203125, 0.0, -86.203125, -57.21875, 91.890625]
  {
    16'b0000000000000000,  // 0.0
    16'b1110100100000111,  // -91.890625
    16'b0000111001001110,  // 57.21875
    16'b0001010110001101,  // 86.203125
    16'b0000000000000000,  // 0.0
    16'b1110101001110011,  // -86.203125
    16'b1111000110110010,  // -57.21875
    16'b0001011011111001   // 91.890625
  },
  // y_im_15 = [0.0, 88.9375, -25.890625, 19.625, 0.0, -19.625, 25.890625, -88.9375]
  {
    16'b0000000000000000,  // 0.0
    16'b0001011000111100,  // 88.9375
    16'b1111100110000111,  // -25.890625
    16'b0000010011101000,  // 19.625
    16'b0000000000000000,  // 0.0
    16'b1111101100011000,  // -19.625
    16'b0000011001111001,  // 25.890625
    16'b1110100111000100   // -88.9375
  },
  // y_im_16 = [0.0, -1.171875, 19.8125, 63.421875, 0.0, -63.421875, -19.8125, 1.171875]
  {
    16'b0000000000000000,  // 0.0
    16'b1111111110110101,  // -1.171875
    16'b0000010011110100,  // 19.8125
    16'b0000111111011011,  // 63.421875
    16'b0000000000000000,  // 0.0
    16'b1111000000100101,  // -63.421875
    16'b1111101100001100,  // -19.8125
    16'b0000000001001011   // 1.171875
  },
  // y_im_17 = [0.0, -31.90625, -14.8125, 97.5, 0.0, -97.5, 14.8125, 31.90625]
  {
    16'b0000000000000000,  // 0.0
    16'b1111100000000110,  // -31.90625
    16'b1111110001001100,  // -14.8125
    16'b0001100001100000,  // 97.5
    16'b0000000000000000,  // 0.0
    16'b1110011110100000,  // -97.5
    16'b0000001110110100,  // 14.8125
    16'b0000011111111010   // 31.90625
  },
  // y_im_18 = [0.0, -38.453125, 131.09375, 43.265625, 0.0, -43.265625, -131.09375, 38.453125]
  {
    16'b0000000000000000,  // 0.0
    16'b1111011001100011,  // -38.453125
    16'b0010000011000110,  // 131.09375
    16'b0000101011010001,  // 43.265625
    16'b0000000000000000,  // 0.0
    16'b1111010100101111,  // -43.265625
    16'b1101111100111010,  // -131.09375
    16'b0000100110011101   // 38.453125
  },
  // y_im_19 = [0.0, 59.375, -27.03125, 78.5, 0.0, -78.5, 27.03125, -59.375]
  {
    16'b0000000000000000,  // 0.0
    16'b0000111011011000,  // 59.375
    16'b1111100100111110,  // -27.03125
    16'b0001001110100000,  // 78.5
    16'b0000000000000000,  // 0.0
    16'b1110110001100000,  // -78.5
    16'b0000011011000010,  // 27.03125
    16'b1111000100101000   // -59.375
  },
  // y_im_20 = [0.0, 2.546875, 39.71875, -31.828125, 0.0, 31.828125, -39.71875, -2.546875]
  {
    16'b0000000000000000,  // 0.0
    16'b0000000010100011,  // 2.546875
    16'b0000100111101110,  // 39.71875
    16'b1111100000001011,  // -31.828125
    16'b0000000000000000,  // 0.0
    16'b0000011111110101,  // 31.828125
    16'b1111011000010010,  // -39.71875
    16'b1111111101011101   // -2.546875
  },
  // y_im_21 = [0.0, -100.140625, -20.453125, -156.453125, 0.0, 156.453125, 20.453125, 100.140625]
  {
    16'b0000000000000000,  // 0.0
    16'b1110011011110111,  // -100.140625
    16'b1111101011100011,  // -20.453125
    16'b1101100011100011,  // -156.453125
    16'b0000000000000000,  // 0.0
    16'b0010011100011101,  // 156.453125
    16'b0000010100011101,  // 20.453125
    16'b0001100100001001   // 100.140625
  },
  // y_im_22 = [0.0, 86.796875, 79.078125, 42.203125, 0.0, -42.203125, -79.078125, -86.796875]
  {
    16'b0000000000000000,  // 0.0
    16'b0001010110110011,  // 86.796875
    16'b0001001111000101,  // 79.078125
    16'b0000101010001101,  // 42.203125
    16'b0000000000000000,  // 0.0
    16'b1111010101110011,  // -42.203125
    16'b1110110000111011,  // -79.078125
    16'b1110101001001101   // -86.796875
  },
  // y_im_23 = [0.0, -23.484375, 137.109375, 103.921875, 0.0, -103.921875, -137.109375, 23.484375]
  {
    16'b0000000000000000,  // 0.0
    16'b1111101000100001,  // -23.484375
    16'b0010001001000111,  // 137.109375
    16'b0001100111111011,  // 103.921875
    16'b0000000000000000,  // 0.0
    16'b1110011000000101,  // -103.921875
    16'b1101110110111001,  // -137.109375
    16'b0000010111011111   // 23.484375
  },
  // y_im_24 = [0.0, -145.0, -52.828125, 104.09375, 0.0, -104.09375, 52.828125, 145.0]
  {
    16'b0000000000000000,  // 0.0
    16'b1101101111000000,  // -145.0
    16'b1111001011001011,  // -52.828125
    16'b0001101000000110,  // 104.09375
    16'b0000000000000000,  // 0.0
    16'b1110010111111010,  // -104.09375
    16'b0000110100110101,  // 52.828125
    16'b0010010001000000   // 145.0
  },
  // y_im_25 = [0.0, 102.125, 82.5, 25.96875, 0.0, -25.96875, -82.5, -102.125]
  {
    16'b0000000000000000,  // 0.0
    16'b0001100110001000,  // 102.125
    16'b0001010010100000,  // 82.5
    16'b0000011001111110,  // 25.96875
    16'b0000000000000000,  // 0.0
    16'b1111100110000010,  // -25.96875
    16'b1110101101100000,  // -82.5
    16'b1110011001111000   // -102.125
  },
  // y_im_26 = [0.0, -0.375, 63.390625, 83.25, 0.0, -83.25, -63.390625, 0.375]
  {
    16'b0000000000000000,  // 0.0
    16'b1111111111101000,  // -0.375
    16'b0000111111011001,  // 63.390625
    16'b0001010011010000,  // 83.25
    16'b0000000000000000,  // 0.0
    16'b1110101100110000,  // -83.25
    16'b1111000000100111,  // -63.390625
    16'b0000000000011000   // 0.375
  },
  // y_im_27 = [0.0, -9.984375, -126.03125, -28.640625, 0.0, 28.640625, 126.03125, 9.984375]
  {
    16'b0000000000000000,  // 0.0
    16'b1111110110000001,  // -9.984375
    16'b1110000001111110,  // -126.03125
    16'b1111100011010111,  // -28.640625
    16'b0000000000000000,  // 0.0
    16'b0000011100101001,  // 28.640625
    16'b0001111110000010,  // 126.03125
    16'b0000001001111111   // 9.984375
  },
  // y_im_28 = [0.0, 39.265625, -63.890625, -151.453125, 0.0, 151.453125, 63.890625, -39.265625]
  {
    16'b0000000000000000,  // 0.0
    16'b0000100111010001,  // 39.265625
    16'b1111000000000111,  // -63.890625
    16'b1101101000100011,  // -151.453125
    16'b0000000000000000,  // 0.0
    16'b0010010111011101,  // 151.453125
    16'b0000111111111001,  // 63.890625
    16'b1111011000101111   // -39.265625
  },
  // y_im_29 = [0.0, -27.046875, -124.734375, 158.921875, 0.0, -158.921875, 124.734375, 27.046875]
  {
    16'b0000000000000000,  // 0.0
    16'b1111100100111101,  // -27.046875
    16'b1110000011010001,  // -124.734375
    16'b0010011110111011,  // 158.921875
    16'b0000000000000000,  // 0.0
    16'b1101100001000101,  // -158.921875
    16'b0001111100101111,  // 124.734375
    16'b0000011011000011   // 27.046875
  },
  // y_im_30 = [0.0, 97.4375, -116.90625, 48.34375, 0.0, -48.34375, 116.90625, -97.4375]
  {
    16'b0000000000000000,  // 0.0
    16'b0001100001011100,  // 97.4375
    16'b1110001011000110,  // -116.90625
    16'b0000110000010110,  // 48.34375
    16'b0000000000000000,  // 0.0
    16'b1111001111101010,  // -48.34375
    16'b0001110100111010,  // 116.90625
    16'b1110011110100100   // -97.4375
  },
  // y_im_31 = [0.0, -57.671875, -32.484375, -110.171875, 0.0, 110.171875, 32.484375, 57.671875]
  {
    16'b0000000000000000,  // 0.0
    16'b1111000110010101,  // -57.671875
    16'b1111011111100001,  // -32.484375
    16'b1110010001110101,  // -110.171875
    16'b0000000000000000,  // 0.0
    16'b0001101110001011,  // 110.171875
    16'b0000100000011111,  // 32.484375
    16'b0000111001101011   // 57.671875
  },
  // y_im_32 = [0.0, 4.625, 88.875, 47.6875, 0.0, -47.6875, -88.875, -4.625]
  {
    16'b0000000000000000,  // 0.0
    16'b0000000100101000,  // 4.625
    16'b0001011000111000,  // 88.875
    16'b0000101111101100,  // 47.6875
    16'b0000000000000000,  // 0.0
    16'b1111010000010100,  // -47.6875
    16'b1110100111001000,  // -88.875
    16'b1111111011011000   // -4.625
  },
  // y_im_33 = [0.0, 15.765625, 2.046875, -69.078125, 0.0, 69.078125, -2.046875, -15.765625]
  {
    16'b0000000000000000,  // 0.0
    16'b0000001111110001,  // 15.765625
    16'b0000000010000011,  // 2.046875
    16'b1110111010111011,  // -69.078125
    16'b0000000000000000,  // 0.0
    16'b0001000101000101,  // 69.078125
    16'b1111111101111101,  // -2.046875
    16'b1111110000001111   // -15.765625
  },
  // y_im_34 = [0.0, 144.65625, 31.578125, 139.28125, 0.0, -139.28125, -31.578125, -144.65625]
  {
    16'b0000000000000000,  // 0.0
    16'b0010010000101010,  // 144.65625
    16'b0000011111100101,  // 31.578125
    16'b0010001011010010,  // 139.28125
    16'b0000000000000000,  // 0.0
    16'b1101110100101110,  // -139.28125
    16'b1111100000011011,  // -31.578125
    16'b1101101111010110   // -144.65625
  },
  // y_im_35 = [0.0, -19.765625, 93.671875, 97.453125, 0.0, -97.453125, -93.671875, 19.765625]
  {
    16'b0000000000000000,  // 0.0
    16'b1111101100001111,  // -19.765625
    16'b0001011101101011,  // 93.671875
    16'b0001100001011101,  // 97.453125
    16'b0000000000000000,  // 0.0
    16'b1110011110100011,  // -97.453125
    16'b1110100010010101,  // -93.671875
    16'b0000010011110001   // 19.765625
  },
  // y_im_36 = [0.0, 85.609375, -37.484375, -105.703125, 0.0, 105.703125, 37.484375, -85.609375]
  {
    16'b0000000000000000,  // 0.0
    16'b0001010101100111,  // 85.609375
    16'b1111011010100001,  // -37.484375
    16'b1110010110010011,  // -105.703125
    16'b0000000000000000,  // 0.0
    16'b0001101001101101,  // 105.703125
    16'b0000100101011111,  // 37.484375
    16'b1110101010011001   // -85.609375
  },
  // y_im_37 = [0.0, 71.6875, 75.65625, 22.5625, 0.0, -22.5625, -75.65625, -71.6875]
  {
    16'b0000000000000000,  // 0.0
    16'b0001000111101100,  // 71.6875
    16'b0001001011101010,  // 75.65625
    16'b0000010110100100,  // 22.5625
    16'b0000000000000000,  // 0.0
    16'b1111101001011100,  // -22.5625
    16'b1110110100010110,  // -75.65625
    16'b1110111000010100   // -71.6875
  },
  // y_im_38 = [0.0, 27.78125, -28.671875, 21.5, 0.0, -21.5, 28.671875, -27.78125]
  {
    16'b0000000000000000,  // 0.0
    16'b0000011011110010,  // 27.78125
    16'b1111100011010101,  // -28.671875
    16'b0000010101100000,  // 21.5
    16'b0000000000000000,  // 0.0
    16'b1111101010100000,  // -21.5
    16'b0000011100101011,  // 28.671875
    16'b1111100100001110   // -27.78125
  },
  // y_im_39 = [0.0, -18.9375, 24.703125, -33.09375, 0.0, 33.09375, -24.703125, 18.9375]
  {
    16'b0000000000000000,  // 0.0
    16'b1111101101000100,  // -18.9375
    16'b0000011000101101,  // 24.703125
    16'b1111011110111010,  // -33.09375
    16'b0000000000000000,  // 0.0
    16'b0000100001000110,  // 33.09375
    16'b1111100111010011,  // -24.703125
    16'b0000010010111100   // 18.9375
  },
  // y_im_40 = [0.0, -43.78125, -59.265625, 83.125, 0.0, -83.125, 59.265625, 43.78125]
  {
    16'b0000000000000000,  // 0.0
    16'b1111010100001110,  // -43.78125
    16'b1111000100101111,  // -59.265625
    16'b0001010011001000,  // 83.125
    16'b0000000000000000,  // 0.0
    16'b1110101100111000,  // -83.125
    16'b0000111011010001,  // 59.265625
    16'b0000101011110010   // 43.78125
  },
  // y_im_41 = [0.0, 37.046875, -57.8125, 22.921875, 0.0, -22.921875, 57.8125, -37.046875]
  {
    16'b0000000000000000,  // 0.0
    16'b0000100101000011,  // 37.046875
    16'b1111000110001100,  // -57.8125
    16'b0000010110111011,  // 22.921875
    16'b0000000000000000,  // 0.0
    16'b1111101001000101,  // -22.921875
    16'b0000111001110100,  // 57.8125
    16'b1111011010111101   // -37.046875
  },
  // y_im_42 = [0.0, 40.609375, 95.65625, -133.765625, 0.0, 133.765625, -95.65625, -40.609375]
  {
    16'b0000000000000000,  // 0.0
    16'b0000101000100111,  // 40.609375
    16'b0001011111101010,  // 95.65625
    16'b1101111010001111,  // -133.765625
    16'b0000000000000000,  // 0.0
    16'b0010000101110001,  // 133.765625
    16'b1110100000010110,  // -95.65625
    16'b1111010111011001   // -40.609375
  },
  // y_im_43 = [0.0, -112.59375, 24.453125, -63.59375, 0.0, 63.59375, -24.453125, 112.59375]
  {
    16'b0000000000000000,  // 0.0
    16'b1110001111011010,  // -112.59375
    16'b0000011000011101,  // 24.453125
    16'b1111000000011010,  // -63.59375
    16'b0000000000000000,  // 0.0
    16'b0000111111100110,  // 63.59375
    16'b1111100111100011,  // -24.453125
    16'b0001110000100110   // 112.59375
  },
  // y_im_44 = [0.0, 45.21875, 26.25, -74.0, 0.0, 74.0, -26.25, -45.21875]
  {
    16'b0000000000000000,  // 0.0
    16'b0000101101001110,  // 45.21875
    16'b0000011010010000,  // 26.25
    16'b1110110110000000,  // -74.0
    16'b0000000000000000,  // 0.0
    16'b0001001010000000,  // 74.0
    16'b1111100101110000,  // -26.25
    16'b1111010010110010   // -45.21875
  },
  // y_im_45 = [0.0, 33.015625, 57.453125, -25.546875, 0.0, 25.546875, -57.453125, -33.015625]
  {
    16'b0000000000000000,  // 0.0
    16'b0000100001000001,  // 33.015625
    16'b0000111001011101,  // 57.453125
    16'b1111100110011101,  // -25.546875
    16'b0000000000000000,  // 0.0
    16'b0000011001100011,  // 25.546875
    16'b1111000110100011,  // -57.453125
    16'b1111011110111111   // -33.015625
  },
  // y_im_46 = [0.0, 6.4375, 9.578125, 103.0, 0.0, -103.0, -9.578125, -6.4375]
  {
    16'b0000000000000000,  // 0.0
    16'b0000000110011100,  // 6.4375
    16'b0000001001100101,  // 9.578125
    16'b0001100111000000,  // 103.0
    16'b0000000000000000,  // 0.0
    16'b1110011001000000,  // -103.0
    16'b1111110110011011,  // -9.578125
    16'b1111111001100100   // -6.4375
  },
  // y_im_47 = [0.0, 49.171875, 167.171875, -29.734375, 0.0, 29.734375, -167.171875, -49.171875]
  {
    16'b0000000000000000,  // 0.0
    16'b0000110001001011,  // 49.171875
    16'b0010100111001011,  // 167.171875
    16'b1111100010010001,  // -29.734375
    16'b0000000000000000,  // 0.0
    16'b0000011101101111,  // 29.734375
    16'b1101011000110101,  // -167.171875
    16'b1111001110110101   // -49.171875
  },
  // y_im_48 = [0.0, -147.546875, 42.71875, 21.609375, 0.0, -21.609375, -42.71875, 147.546875]
  {
    16'b0000000000000000,  // 0.0
    16'b1101101100011101,  // -147.546875
    16'b0000101010101110,  // 42.71875
    16'b0000010101100111,  // 21.609375
    16'b0000000000000000,  // 0.0
    16'b1111101010011001,  // -21.609375
    16'b1111010101010010,  // -42.71875
    16'b0010010011100011   // 147.546875
  },
  // y_im_49 = [0.0, -29.484375, -130.671875, 2.203125, 0.0, -2.203125, 130.671875, 29.484375]
  {
    16'b0000000000000000,  // 0.0
    16'b1111100010100001,  // -29.484375
    16'b1101111101010101,  // -130.671875
    16'b0000000010001101,  // 2.203125
    16'b0000000000000000,  // 0.0
    16'b1111111101110011,  // -2.203125
    16'b0010000010101011,  // 130.671875
    16'b0000011101011111   // 29.484375
  },
  // y_im_50 = [0.0, -67.421875, 17.15625, 15.765625, 0.0, -15.765625, -17.15625, 67.421875]
  {
    16'b0000000000000000,  // 0.0
    16'b1110111100100101,  // -67.421875
    16'b0000010001001010,  // 17.15625
    16'b0000001111110001,  // 15.765625
    16'b0000000000000000,  // 0.0
    16'b1111110000001111,  // -15.765625
    16'b1111101110110110,  // -17.15625
    16'b0001000011011011   // 67.421875
  },
  // y_im_51 = [0.0, 87.40625, -60.265625, 124.03125, 0.0, -124.03125, 60.265625, -87.40625]
  {
    16'b0000000000000000,  // 0.0
    16'b0001010111011010,  // 87.40625
    16'b1111000011101111,  // -60.265625
    16'b0001111100000010,  // 124.03125
    16'b0000000000000000,  // 0.0
    16'b1110000011111110,  // -124.03125
    16'b0000111100010001,  // 60.265625
    16'b1110101000100110   // -87.40625
  },
  // y_im_52 = [0.0, 38.5, -80.625, -78.46875, 0.0, 78.46875, 80.625, -38.5]
  {
    16'b0000000000000000,  // 0.0
    16'b0000100110100000,  // 38.5
    16'b1110101111011000,  // -80.625
    16'b1110110001100010,  // -78.46875
    16'b0000000000000000,  // 0.0
    16'b0001001110011110,  // 78.46875
    16'b0001010000101000,  // 80.625
    16'b1111011001100000   // -38.5
  },
  // y_im_53 = [0.0, 45.5625, -54.71875, -87.6875, 0.0, 87.6875, 54.71875, -45.5625]
  {
    16'b0000000000000000,  // 0.0
    16'b0000101101100100,  // 45.5625
    16'b1111001001010010,  // -54.71875
    16'b1110101000010100,  // -87.6875
    16'b0000000000000000,  // 0.0
    16'b0001010111101100,  // 87.6875
    16'b0000110110101110,  // 54.71875
    16'b1111010010011100   // -45.5625
  },
  // y_im_54 = [0.0, -64.84375, -100.65625, 108.0625, 0.0, -108.0625, 100.65625, 64.84375]
  {
    16'b0000000000000000,  // 0.0
    16'b1110111111001010,  // -64.84375
    16'b1110011011010110,  // -100.65625
    16'b0001101100000100,  // 108.0625
    16'b0000000000000000,  // 0.0
    16'b1110010011111100,  // -108.0625
    16'b0001100100101010,  // 100.65625
    16'b0001000000110110   // 64.84375
  },
  // y_im_55 = [0.0, 13.890625, -184.6875, -21.640625, 0.0, 21.640625, 184.6875, -13.890625]
  {
    16'b0000000000000000,  // 0.0
    16'b0000001101111001,  // 13.890625
    16'b1101000111010100,  // -184.6875
    16'b1111101010010111,  // -21.640625
    16'b0000000000000000,  // 0.0
    16'b0000010101101001,  // 21.640625
    16'b0010111000101100,  // 184.6875
    16'b1111110010000111   // -13.890625
  },
  // y_im_56 = [0.0, -6.796875, -24.875, 18.953125, 0.0, -18.953125, 24.875, 6.796875]
  {
    16'b0000000000000000,  // 0.0
    16'b1111111001001101,  // -6.796875
    16'b1111100111001000,  // -24.875
    16'b0000010010111101,  // 18.953125
    16'b0000000000000000,  // 0.0
    16'b1111101101000011,  // -18.953125
    16'b0000011000111000,  // 24.875
    16'b0000000110110011   // 6.796875
  },
  // y_im_57 = [0.0, -48.015625, 168.078125, 77.671875, 0.0, -77.671875, -168.078125, 48.015625]
  {
    16'b0000000000000000,  // 0.0
    16'b1111001111111111,  // -48.015625
    16'b0010101000000101,  // 168.078125
    16'b0001001101101011,  // 77.671875
    16'b0000000000000000,  // 0.0
    16'b1110110010010101,  // -77.671875
    16'b1101010111111011,  // -168.078125
    16'b0000110000000001   // 48.015625
  },
  // y_im_58 = [0.0, -52.078125, -35.078125, 47.140625, 0.0, -47.140625, 35.078125, 52.078125]
  {
    16'b0000000000000000,  // 0.0
    16'b1111001011111011,  // -52.078125
    16'b1111011100111011,  // -35.078125
    16'b0000101111001001,  // 47.140625
    16'b0000000000000000,  // 0.0
    16'b1111010000110111,  // -47.140625
    16'b0000100011000101,  // 35.078125
    16'b0000110100000101   // 52.078125
  },
  // y_im_59 = [0.0, 79.1875, -51.921875, 68.03125, 0.0, -68.03125, 51.921875, -79.1875]
  {
    16'b0000000000000000,  // 0.0
    16'b0001001111001100,  // 79.1875
    16'b1111001100000101,  // -51.921875
    16'b0001000100000010,  // 68.03125
    16'b0000000000000000,  // 0.0
    16'b1110111011111110,  // -68.03125
    16'b0000110011111011,  // 51.921875
    16'b1110110000110100   // -79.1875
  },
  // y_im_60 = [0.0, -119.5625, 27.796875, 91.125, 0.0, -91.125, -27.796875, 119.5625]
  {
    16'b0000000000000000,  // 0.0
    16'b1110001000011100,  // -119.5625
    16'b0000011011110011,  // 27.796875
    16'b0001011011001000,  // 91.125
    16'b0000000000000000,  // 0.0
    16'b1110100100111000,  // -91.125
    16'b1111100100001101,  // -27.796875
    16'b0001110111100100   // 119.5625
  },
  // y_im_61 = [0.0, -57.859375, 144.96875, 10.796875, 0.0, -10.796875, -144.96875, 57.859375]
  {
    16'b0000000000000000,  // 0.0
    16'b1111000110001001,  // -57.859375
    16'b0010010000111110,  // 144.96875
    16'b0000001010110011,  // 10.796875
    16'b0000000000000000,  // 0.0
    16'b1111110101001101,  // -10.796875
    16'b1101101111000010,  // -144.96875
    16'b0000111001110111   // 57.859375
  },
  // y_im_62 = [0.0, 19.046875, -69.109375, 52.953125, 0.0, -52.953125, 69.109375, -19.046875]
  {
    16'b0000000000000000,  // 0.0
    16'b0000010011000011,  // 19.046875
    16'b1110111010111001,  // -69.109375
    16'b0000110100111101,  // 52.953125
    16'b0000000000000000,  // 0.0
    16'b1111001011000011,  // -52.953125
    16'b0001000101000111,  // 69.109375
    16'b1111101100111101   // -19.046875
  },
  // y_im_63 = [0.0, -171.421875, 22.671875, -43.046875, 0.0, 43.046875, -22.671875, 171.421875]
  {
    16'b0000000000000000,  // 0.0
    16'b1101010100100101,  // -171.421875
    16'b0000010110101011,  // 22.671875
    16'b1111010100111101,  // -43.046875
    16'b0000000000000000,  // 0.0
    16'b0000101011000011,  // 43.046875
    16'b1111101001010101,  // -22.671875
    16'b0010101011011011   // 171.421875
  }
};

endpackage