////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2020 Fredrik Åkerlund
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <https://www.gnu.org/licenses/>.
//
// Description:
//
////////////////////////////////////////////////////////////////////////////////

`ifndef CORDIC_AXI4S_TYPES_PKG
`define CORDIC_AXI4S_TYPES_PKG

package cordic_axi4s_types_pkg;

  typedef enum {
    CORDIC_SINE_E,
    CORDIC_COSINE_E,
    CORDIC_SINE_COSINE_E
  } cordic_request_t;

endpackage

`endif
