////////////////////////////////////////////////////////////////////////////////
//
// Copyright 2020 Fredrik Åkerlund
//
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either
// version 2.1 of the License, or (at your option) any later version.
//
// This library is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public
// License along with this library; if not, write to the Free Software
// Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA 02110-1301, USA
//
// Description:
//
////////////////////////////////////////////////////////////////////////////////

`ifndef CORDIC_ATAN_RADIAN_TABLE_PKG
`define CORDIC_ATAN_RADIAN_TABLE_PKG

package cordic_atan_radian_table_pkg;

  // Positive values of n/4*pi in fixed point representation
  localparam logic signed [53 : 0] pi_2_4_pos_n4_q50 = 54'b000110010010000111111011010101000100010000101101000110; // 90  deg  |  1.570796326795 rad | pi/2
  localparam logic signed [53 : 0] pi_4_4_pos_n4_q50 = 54'b001100100100001111110110101010001000100001011010001100; // 180 deg  |  3.141592653590 rad | pi
  localparam logic signed [53 : 0] pi_6_4_pos_n4_q50 = 54'b010010110110010111110001111111001100110010000111010010; // 270 deg  |  4.712388980385 rad | pi*6/4
  localparam logic signed [53 : 0] pi_8_4_pos_n4_q50 = 54'b011001001000011111101101010100010001000010110100011000; // 360 deg  |  6.283185307180 rad | pi*2

  // Negative values of n/4*pi in fixed point representation
  localparam logic signed [53 : 0] pi_2_4_neg_n4_q50 = 54'b111001101101111000000100101010111011101111010010111010; // -90  deg | -1.570796326795 rad | -pi/2
  localparam logic signed [53 : 0] pi_4_4_neg_n4_q50 = 54'b110011011011110000001001010101110111011110100101110100; // -180 deg | -3.141592653590 rad | -pi
  localparam logic signed [53 : 0] pi_6_4_neg_n4_q50 = 54'b101101001001101000001110000000110011001101111000101110; // -270 deg | -4.712388980385 rad | -pi*6/4

  // This table contains a fixed point representation in radians of the rotating
  // theta vector in the CORDIC algorithm.
  localparam logic signed [63 : 0] atan_radian_table_32stage_n4q60 [31] = {
    64'b0000110010010000111111011010101000100010000101101000110000000000, // atan(2^-0)  -> 45.000000000 degrees -> 0.785398163 radians
    64'b0000011101101011000110011100000101011000011011101101001111000000, // atan(2^-1)  -> 26.565051177 degrees -> 0.463647609 radians
    64'b0000001111101011011011101011111100100101100100000001101110100000, // atan(2^-2)  -> 14.036243468 degrees -> 0.244978663 radians
    64'b0000000111111101010110111010100110101010110000101111011011100000, // atan(2^-3)  ->  7.125016349 degrees -> 0.124354995 radians
    64'b0000000011111111101010101101110110111001011001111110111101010000, // atan(2^-4)  ->  3.576334375 degrees -> 0.062418810 radians
    64'b0000000001111111111101010101011011101110101001011101100010010100, // atan(2^-5)  ->  1.789910608 degrees -> 0.031239833 radians
    64'b0000000000111111111111101010101010110111011101101110010100110110, // atan(2^-6)  ->  0.895173710 degrees -> 0.015623729 radians
    64'b0000000000011111111111111101010101010101101110111011101010010111, // atan(2^-7)  ->  0.447614171 degrees -> 0.007812341 radians
    64'b0000000000001111111111111111101010101010101011011101110111011011, // atan(2^-8)  ->  0.223810500 degrees -> 0.003906230 radians
    64'b0000000000000111111111111111111101010101010101010110111011101111, // atan(2^-9)  ->  0.111905677 degrees -> 0.001953123 radians
    64'b0000000000000011111111111111111111101010101010101010101101110111, // atan(2^-10) ->  0.055952892 degrees -> 0.000976562 radians
    64'b0000000000000001111111111111111111111101010101010101010101011011, // atan(2^-11) ->  0.027976453 degrees -> 0.000488281 radians
    64'b0000000000000000111111111111111111111111101010101010101010101010, // atan(2^-12) ->  0.013988227 degrees -> 0.000244141 radians
    64'b0000000000000000011111111111111111111111111101010101010101010101, // atan(2^-13) ->  0.006994114 degrees -> 0.000122070 radians
    64'b0000000000000000001111111111111111111111111111101010101010101010, // atan(2^-14) ->  0.003497057 degrees -> 0.000061035 radians
    64'b0000000000000000000111111111111111111111111111111101010101010101, // atan(2^-15) ->  0.001748528 degrees -> 0.000030518 radians
    64'b0000000000000000000011111111111111111111111111111111101010101010, // atan(2^-16) ->  0.000874264 degrees -> 0.000015259 radians
    64'b0000000000000000000001111111111111111111111111111111111101010101, // atan(2^-17) ->  0.000437132 degrees -> 0.000007629 radians
    64'b0000000000000000000000111111111111111111111111111111111111101010, // atan(2^-18) ->  0.000218566 degrees -> 0.000003815 radians
    64'b0000000000000000000000011111111111111111111111111111111111111101, // atan(2^-19) ->  0.000109283 degrees -> 0.000001907 radians
    64'b0000000000000000000000001111111111111111111111111111111111111111, // atan(2^-20) ->  0.000054642 degrees -> 0.000000954 radians
    64'b0000000000000000000000000111111111111111111111111111111111111111, // atan(2^-21) ->  0.000027321 degrees -> 0.000000477 radians
    64'b0000000000000000000000000011111111111111111111111111111111111111, // atan(2^-22) ->  0.000013660 degrees -> 0.000000238 radians
    64'b0000000000000000000000000001111111111111111111111111111111111111, // atan(2^-23) ->  0.000006830 degrees -> 0.000000119 radians
    64'b0000000000000000000000000000111111111111111111111111111111111111, // atan(2^-24) ->  0.000003415 degrees -> 0.000000060 radians
    64'b0000000000000000000000000000011111111111111111111111111111111111, // atan(2^-25) ->  0.000001708 degrees -> 0.000000030 radians
    64'b0000000000000000000000000000001111111111111111111111111111111111, // atan(2^-26) ->  0.000000854 degrees -> 0.000000015 radians
    64'b0000000000000000000000000000001000000000000000000000000000000000, // atan(2^-27) ->  0.000000427 degrees -> 0.000000007 radians
    64'b0000000000000000000000000000000100000000000000000000000000000000, // atan(2^-28) ->  0.000000213 degrees -> 0.000000004 radians
    64'b0000000000000000000000000000000010000000000000000000000000000000, // atan(2^-29) ->  0.000000107 degrees -> 0.000000002 radians
    64'b0000000000000000000000000000000001000000000000000000000000000000  // atan(2^-30) ->  0.000000053 degrees -> 0.000000001 radians
  };

  // This table contains a fixed point representation of the gain that is
  // inherent from the CORDIC algorithm. Depending on how many stages that
  // are used, one of these vectors shall be assinged as the input X vector.
  localparam logic signed [63 : 0] gain_table_32stage_n4q60 [31] = {
    64'b0000101101010000010011110011001100111111100111011110011000000000, // -> 0.707106781187 (Gain for 1  stages = 1.414213562373)
    64'b0000101000011110100010011011000100100100001001001000011110000000, // -> 0.632455532034 (Gain for 2  stages = 1.581138830084)
    64'b0000100111010001001100001101110100110110101111010001101100000000, // -> 0.613571991078 (Gain for 3  stages = 1.629800601301)
    64'b0000100110111101110010001010000011101111010110011111111100000000, // -> 0.608833912518 (Gain for 4  stages = 1.642484065752)
    64'b0000100110111000111011010110000011000001011101110111101010000000, // -> 0.607648256256 (Gain for 5  stages = 1.645688915757)
    64'b0000100110110111101101100111110101011110110010110000111110000000, // -> 0.607351770141 (Gain for 6  stages = 1.646492278712)
    64'b0000100110110111011010001100001101001111100100111111010010000000, // -> 0.607277644094 (Gain for 7  stages = 1.646693254274)
    64'b0000100110110111010101010101010010111000010110010000100000000000, // -> 0.607259112299 (Gain for 8  stages = 1.646743506597)
    64'b0000100110110111010100000111100100010001010100110110100010000000, // -> 0.607254479333 (Gain for 9  stages = 1.646756070205)
    64'b0000100110110111010011110100001000100111011111101001001000000000, // -> 0.607253321090 (Gain for 10 stages = 1.646759211140)
    64'b0000100110110111010011101111010001101101000010000010010110000000, // -> 0.607253031529 (Gain for 11 stages = 1.646759996376)
    64'b0000100110110111010011101110000011111110011010100111011100000000, // -> 0.607252959139 (Gain for 12 stages = 1.646760192685)
    64'b0000100110110111010011101101110000100010110000110000101010000000, // -> 0.607252941041 (Gain for 13 stages = 1.646760241762)
    64'b0000100110110111010011101101101011101011110110010010111100000000, // -> 0.607252936517 (Gain for 14 stages = 1.646760254031)
    64'b0000100110110111010011101101101010011110000111101011100000000000, // -> 0.607252935386 (Gain for 15 stages = 1.646760257099)
    64'b0000100110110111010011101101101010001010101100000001101010000000, // -> 0.607252935103 (Gain for 16 stages = 1.646760257865)
    64'b0000100110110111010011101101101010000101110101000111001010000000, // -> 0.607252935032 (Gain for 17 stages = 1.646760258057)
    64'b0000100110110111010011101101101010000100100111011000100100000000, // -> 0.607252935015 (Gain for 18 stages = 1.646760258105)
    64'b0000100110110111010011101101101010000100010011111100111010000000, // -> 0.607252935010 (Gain for 19 stages = 1.646760258117)
    64'b0000100110110111010011101101101010000100001111000110000000000000, // -> 0.607252935009 (Gain for 20 stages = 1.646760258120)
    64'b0000100110110111010011101101101010000100001101111000010000000000, // -> 0.607252935009 (Gain for 21 stages = 1.646760258121)
    64'b0000100110110111010011101101101010000100001101100100110110000000, // -> 0.607252935009 (Gain for 22 stages = 1.646760258121)
    64'b0000100110110111010011101101101010000100001101011111111110000000, // -> 0.607252935009 (Gain for 23 stages = 1.646760258121)
    64'b0000100110110111010011101101101010000100001101011110110000000000, // -> 0.607252935009 (Gain for 24 stages = 1.646760258121)
    64'b0000100110110111010011101101101010000100001101011110011100000000, // -> 0.607252935009 (Gain for 25 stages = 1.646760258121)
    64'b0000100110110111010011101101101010000100001101011110011000000000, // -> 0.607252935009 (Gain for 26 stages = 1.646760258121)
    64'b0000100110110111010011101101101010000100001101011110011000000000, // -> 0.607252935009 (Gain for 27 stages = 1.646760258121)
    64'b0000100110110111010011101101101010000100001101011110011000000000, // -> 0.607252935009 (Gain for 28 stages = 1.646760258121)
    64'b0000100110110111010011101101101010000100001101011110011000000000, // -> 0.607252935009 (Gain for 29 stages = 1.646760258121)
    64'b0000100110110111010011101101101010000100001101011110011000000000, // -> 0.607252935009 (Gain for 30 stages = 1.646760258121)
    64'b0000100110110111010011101101101010000100001101011110011000000000  // -> 0.607252935009 (Gain for 31 stages = 1.646760258121)
  };

endpackage

`endif
