////////////////////////////////////////////////////////////////////////////////
//
// Copyright 2020 Fredrik Åkerlund
//
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either
// version 2.1 of the License, or (at your option) any later version.
//
// This library is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public
// License along with this library; if not, write to the Free Software
// Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA 02110-1301, USA
//
// Description:
//
////////////////////////////////////////////////////////////////////////////////

interface vip_apb3_if #(
    parameter vip_apb3_cfg_t cfg = '{default: '0}
  )(
    input clk,
    input rst_n
  );

  logic [cfg.APB_ADDR_WIDTH_P-1 : 0] paddr;
  logic                              psel;
  logic                              penable;
  logic                              pwrite;
  logic [cfg.APB_DATA_WIDTH_P-1 : 0] pwdata;
  logic                              pready;
  logic [cfg.APB_DATA_WIDTH_P-1 : 0] prdata;
  logic                              pslverr;

endinterface
