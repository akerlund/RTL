package gf_ref_pkg;

localparam int M_C        = 8;
localparam int P_ORDER_C  = 256;
localparam int REF_SIZE_C = 16;

localparam logic [M_C-1 : 0] GF_ADD_C [REF_SIZE_C] [3] = '{
  '{158,150,8},
  '{208,16,192},
  '{96,25,121},
  '{36,163,135},
  '{121,230,159},
  '{252,33,221},
  '{47,24,55},
  '{17,14,31},
  '{92,204,144},
  '{234,77,167},
  '{21,75,94},
  '{24,76,84},
  '{1,212,213},
  '{220,2,222},
  '{59,140,183},
  '{189,55,138}
};

localparam logic [M_C-1 : 0] GF_MUL_C [REF_SIZE_C] [3] = '{
  '{147,26,58},
  '{81,204,115},
  '{57,65,251},
  '{213,137,158},
  '{236,221,39},
  '{101,31,47},
  '{54,3,90},
  '{3,133,148},
  '{88,104,242},
  '{149,209,136},
  '{227,31,116},
  '{42,170,244},
  '{212,132,68},
  '{127,171,210},
  '{96,157,106},
  '{69,87,12}
};

localparam logic [M_C-1 : 0] GF_DIV_C [REF_SIZE_C] [3] = '{
  '{9,150,97},
  '{213,179,97},
  '{10,111,97},
  '{0,198,97},
  '{74,240,97},
  '{94,181,97},
  '{53,176,97},
  '{8,176,97},
  '{160,112,97},
  '{125,110,97},
  '{4,141,97},
  '{218,100,97},
  '{2,67,97},
  '{148,75,97},
  '{153,88,97},
  '{105,233,97}
};

endpackage
