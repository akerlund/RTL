package gf_ref_pkg;

  localparam int M_C        = 8;
  localparam int REF_SIZE_C = 64;

  localparam logic [M_C-1 : 0] GF_ADD_C [REF_SIZE_C] [3] = '{
    '{232,46,198},
    '{122,57,67},
    '{51,214,229},
    '{1,82,83},
    '{29,127,98},
    '{25,16,9},
    '{203,180,127},
    '{115,101,22},
    '{129,243,114},
    '{251,255,4},
    '{91,150,205},
    '{55,148,163},
    '{251,186,65},
    '{117,0,117},
    '{100,87,51},
    '{18,85,71},
    '{185,211,106},
    '{189,79,242},
    '{160,145,49},
    '{182,196,114},
    '{132,96,228},
    '{242,125,143},
    '{127,136,247},
    '{64,250,186},
    '{18,70,84},
    '{244,134,114},
    '{165,247,82},
    '{69,209,148},
    '{222,250,36},
    '{209,250,43},
    '{78,84,26},
    '{169,138,35},
    '{76,236,160},
    '{179,202,121},
    '{56,249,193},
    '{210,45,255},
    '{254,153,103},
    '{228,220,56},
    '{47,36,11},
    '{6,87,81},
    '{152,196,92},
    '{68,9,77},
    '{178,29,175},
    '{224,31,255},
    '{238,74,164},
    '{0,27,27},
    '{191,26,165},
    '{30,163,189},
    '{142,37,171},
    '{127,57,70},
    '{226,221,63},
    '{1,248,249},
    '{75,23,92},
    '{241,59,202},
    '{44,106,70},
    '{154,135,29},
    '{232,50,218},
    '{45,245,216},
    '{204,136,68},
    '{221,20,201},
    '{148,149,1},
    '{69,58,127},
    '{185,14,183},
    '{5,110,107}
  };

  localparam logic [M_C-1 : 0] GF_MUL_C [REF_SIZE_C] [3] = '{
    '{228,214,88},
    '{111,74,67},
    '{202,119,248},
    '{220,60,58},
    '{84,229,186},
    '{153,92,14},
    '{139,249,200},
    '{50,244,229},
    '{26,165,148},
    '{122,43,130},
    '{206,251,223},
    '{79,62,108},
    '{205,177,67},
    '{17,151,18},
    '{248,86,253},
    '{221,244,75},
    '{51,222,220},
    '{80,120,184},
    '{7,38,242},
    '{203,237,67},
    '{133,6,57},
    '{252,120,207},
    '{95,150,250},
    '{70,140,175},
    '{223,225,75},
    '{187,125,188},
    '{85,217,207},
    '{143,53,161},
    '{19,151,33},
    '{138,232,243},
    '{201,204,85},
    '{236,91,249},
    '{151,87,105},
    '{187,202,228},
    '{135,140,222},
    '{207,190,93},
    '{10,203,157},
    '{102,87,185},
    '{12,220,249},
    '{83,203,220},
    '{180,125,29},
    '{198,108,115},
    '{58,189,199},
    '{15,177,209},
    '{109,169,135},
    '{47,186,102},
    '{135,175,103},
    '{163,8,113},
    '{232,223,34},
    '{245,213,109},
    '{120,214,99},
    '{15,187,183},
    '{44,107,47},
    '{84,204,38},
    '{219,165,103},
    '{3,187,208},
    '{19,8,152},
    '{182,107,219},
    '{1,218,218},
    '{60,75,2},
    '{17,224,70},
    '{29,143,157},
    '{84,91,235},
    '{223,105,82}
  };

  localparam logic [M_C-1 : 0] GF_DIV_C [REF_SIZE_C] [3] = '{
    '{236,109,250},
    '{19,67,179},
    '{157,46,213},
    '{114,34,80},
    '{185,245,107},
    '{53,78,32},
    '{224,38,165},
    '{145,233,255},
    '{46,206,90},
    '{90,208,63},
    '{92,179,239},
    '{113,71,217},
    '{16,250,38},
    '{29,126,217},
    '{175,24,47},
    '{102,35,240},
    '{150,108,55},
    '{234,3,173},
    '{233,45,144},
    '{91,135,240},
    '{164,225,185},
    '{157,201,58},
    '{121,67,62},
    '{38,179,134},
    '{55,56,22},
    '{141,69,245},
    '{192,135,45},
    '{154,185,177},
    '{73,175,160},
    '{161,49,158},
    '{199,137,238},
    '{194,203,177},
    '{107,241,145},
    '{170,48,236},
    '{103,193,190},
    '{70,35,2},
    '{116,45,131},
    '{188,159,3},
    '{206,26,64},
    '{224,35,228},
    '{148,64,157},
    '{218,66,108},
    '{182,229,75},
    '{175,28,73},
    '{102,166,241},
    '{184,96,68},
    '{157,244,186},
    '{16,21,199},
    '{93,29,70},
    '{28,82,20},
    '{142,205,176},
    '{132,59,180},
    '{164,204,234},
    '{128,64,2},
    '{3,177,50},
    '{120,100,33},
    '{118,157,225},
    '{51,123,81},
    '{183,55,61},
    '{200,167,207},
    '{158,222,15},
    '{14,241,3},
    '{35,253,138},
    '{149,67,177}
  };

  endpackage
