////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2020 Fredrik Åkerlund
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <https://www.gnu.org/licenses/>.
//
// Description:
//
////////////////////////////////////////////////////////////////////////////////

class tc_awa_basic_write extends awa_base_test;

  awa_write_vseq #(vip_axi4_cfg) awa_write_all;

  `uvm_component_utils(tc_awa_basic_write)



  function new(string name = "tc_awa_basic_write", uvm_component parent = null);

    super.new(name, parent);

    // Memory Agent configuration
    use_response_channel         = 1;
    wready_back_pressure_enabled = 1;

    // Memory Agent configuration
    memory_depth = 16;

  endfunction



  function void build_phase(uvm_phase phase);

    super.build_phase(phase);

  endfunction



  task run_phase(uvm_phase phase);

    super.run_phase(phase);
    phase.raise_objection(this);

    awa_write_all = new();
    awa_write_all.max_awaddr              = 2**memory_depth-1;
    awa_write_all.nr_of_bursts            = 5000;
    awa_write_all.max_idle_between_bursts = 512;
    awa_write_all.start(v_sqr);

    phase.drop_objection(this);

  endtask

endclass
