////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2020 Fredrik Åkerlund
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <https://www.gnu.org/licenses/>.
//
// Description:
//
////////////////////////////////////////////////////////////////////////////////

`ifndef CORDIC_TEST_ANGLES_PKG
`define CORDIC_TEST_ANGLES_PKG

package cordic_test_angles_pkg;

  logic [31 : 0] neg_radians [360] = {
    32'b00000000000000000000000000000000,
    32'b11111111101110001000001011100110,
    32'b11111111011100010000010111001011,
    32'b11111111001010011000100010110001,
    32'b11111110111000100000101110010110,
    32'b11111110100110101000111001111100,
    32'b11111110010100110001000101100001,
    32'b11111110000010111001010001000111,
    32'b11111101110001000001011100101100,
    32'b11111101011111001001101000010010,
    32'b11111101001101010001110011110111,
    32'b11111100111011011001111111011101,
    32'b11111100101001100010001011000010,
    32'b11111100010111101010010110101000,
    32'b11111100000101110010100010001101,
    32'b11111011110011111010101101110010,
    32'b11111011100010000010111001011000,
    32'b11111011010000001011000100111101,
    32'b11111010111110010011010000100011,
    32'b11111010101100011011011100001000,
    32'b11111010011010100011100111101110,
    32'b11111010001000101011110011010011,
    32'b11111001110110110011111110111001,
    32'b11111001100100111100001010011110,
    32'b11111001010011000100010110000100,
    32'b11111001000001001100100001101001,
    32'b11111000101111010100101101001111,
    32'b11111000011101011100111000110100,
    32'b11111000001011100101000100011001,
    32'b11110111111001101101001111111111,
    32'b11110111100111110101011011100100,
    32'b11110111010101111101100111001010,
    32'b11110111000100000101110010101111,
    32'b11110110110010001101111110010101,
    32'b11110110100000010110001001111010,
    32'b11110110001110011110010101100000,
    32'b11110101111100100110100001000101,
    32'b11110101101010101110101100101011,
    32'b11110101011000110110111000010000,
    32'b11110101000110111111000011110110,
    32'b11110100110101000111001111011011,
    32'b11110100100011001111011011000001,
    32'b11110100010001010111100110100110,
    32'b11110011111111011111110010001011,
    32'b11110011101101100111111101110001,
    32'b11110011011011110000001001010110,
    32'b11110011001001111000010100111100,
    32'b11110010111000000000100000100001,
    32'b11110010100110001000101100000111,
    32'b11110010010100010000110111101100,
    32'b11110010000010011001000011010010,
    32'b11110001110000100001001110110111,
    32'b11110001011110101001011010011101,
    32'b11110001001100110001100110000010,
    32'b11110000111010111001110001101000,
    32'b11110000101001000001111101001101,
    32'b11110000010111001010001000110010,
    32'b11110000000101010010010100011000,
    32'b11101111110011011010011111111101,
    32'b11101111100001100010101011100011,
    32'b11101111001111101010110111001000,
    32'b11101110111101110011000010101110,
    32'b11101110101011111011001110010011,
    32'b11101110011010000011011001111001,
    32'b11101110001000001011100101011110,
    32'b11101101110110010011110001000100,
    32'b11101101100100011011111100101001,
    32'b11101101010010100100001000001111,
    32'b11101101000000101100010011110100,
    32'b11101100101110110100011111011001,
    32'b11101100011100111100101010111111,
    32'b11101100001011000100110110100100,
    32'b11101011111001001101000010001010,
    32'b11101011100111010101001101101111,
    32'b11101011010101011101011001010101,
    32'b11101011000011100101100100111010,
    32'b11101010110001101101110000100000,
    32'b11101010011111110101111100000101,
    32'b11101010001101111110000111101011,
    32'b11101001111100000110010011010000,
    32'b11101001101010001110011110110110,
    32'b11101001011000010110101010011011,
    32'b11101001000110011110110110000001,
    32'b11101000110100100111000001100110,
    32'b11101000100010101111001101001011,
    32'b11101000010000110111011000110001,
    32'b11100111111110111111100100010110,
    32'b11100111101101000111101111111100,
    32'b11100111011011001111111011100001,
    32'b11100111001001011000000111000111,
    32'b11100110110111100000010010101100,
    32'b11100110100101101000011110010010,
    32'b11100110010011110000101001110111,
    32'b11100110000001111000110101011101,
    32'b11100101110000000001000001000010,
    32'b11100101011110001001001100101000,
    32'b11100101001100010001011000001101,
    32'b11100100111010011001100011110010,
    32'b11100100101000100001101111011000,
    32'b11100100010110101001111010111101,
    32'b11100100000100110010000110100011,
    32'b11100011110010111010010010001000,
    32'b11100011100001000010011101101110,
    32'b11100011001111001010101001010011,
    32'b11100010111101010010110100111001,
    32'b11100010101011011011000000011110,
    32'b11100010011001100011001100000100,
    32'b11100010000111101011010111101001,
    32'b11100001110101110011100011001111,
    32'b11100001100011111011101110110100,
    32'b11100001010010000011111010011010,
    32'b11100001000000001100000101111111,
    32'b11100000101110010100010001100100,
    32'b11100000011100011100011101001010,
    32'b11100000001010100100101000101111,
    32'b11011111111000101100110100010101,
    32'b11011111100110110100111111111010,
    32'b11011111010100111101001011100000,
    32'b11011111000011000101010111000101,
    32'b11011110110001001101100010101011,
    32'b11011110011111010101101110010000,
    32'b11011110001101011101111001110110,
    32'b11011101111011100110000101011011,
    32'b11011101101001101110010001000001,
    32'b11011101010111110110011100100110,
    32'b11011101000101111110101000001011,
    32'b11011100110100000110110011110001,
    32'b11011100100010001110111111010110,
    32'b11011100010000010111001010111100,
    32'b11011011111110011111010110100001,
    32'b11011011101100100111100010000111,
    32'b11011011011010101111101101101100,
    32'b11011011001000110111111001010010,
    32'b11011010110111000000000100110111,
    32'b11011010100101001000010000011101,
    32'b11011010010011010000011100000010,
    32'b11011010000001011000100111101000,
    32'b11011001101111100000110011001101,
    32'b11011001011101101000111110110010,
    32'b11011001001011110001001010011000,
    32'b11011000111001111001010101111101,
    32'b11011000101000000001100001100011,
    32'b11011000010110001001101101001000,
    32'b11011000000100010001111000101110,
    32'b11010111110010011010000100010011,
    32'b11010111100000100010001111111001,
    32'b11010111001110101010011011011110,
    32'b11010110111100110010100111000100,
    32'b11010110101010111010110010101001,
    32'b11010110011001000010111110001111,
    32'b11010110000111001011001001110100,
    32'b11010101110101010011010101011010,
    32'b11010101100011011011100000111111,
    32'b11010101010001100011101100100100,
    32'b11010100111111101011111000001010,
    32'b11010100101101110100000011101111,
    32'b11010100011011111100001111010101,
    32'b11010100001010000100011010111010,
    32'b11010011111000001100100110100000,
    32'b11010011100110010100110010000101,
    32'b11010011010100011100111101101011,
    32'b11010011000010100101001001010000,
    32'b11010010110000101101010100110110,
    32'b11010010011110110101100000011011,
    32'b11010010001100111101101100000001,
    32'b11010001111011000101110111100110,
    32'b11010001101001001110000011001011,
    32'b11010001010111010110001110110001,
    32'b11010001000101011110011010010110,
    32'b11010000110011100110100101111100,
    32'b11010000100001101110110001100001,
    32'b11010000001111110110111101000111,
    32'b11001111111101111111001000101100,
    32'b11001111101100000111010100010010,
    32'b11001111011010001111011111110111,
    32'b11001111001000010111101011011101,
    32'b11001110110110011111110111000010,
    32'b11001110100100101000000010101000,
    32'b11001110010010110000001110001101,
    32'b11001110000000111000011001110011,
    32'b11001101101111000000100101011000,
    32'b11001101011101001000110000111101,
    32'b11001101001011010000111100100011,
    32'b11001100111001011001001000001000,
    32'b11001100100111100001010011101110,
    32'b11001100010101101001011111010011,
    32'b11001100000011110001101010111001,
    32'b11001011110001111001110110011110,
    32'b11001011100000000010000010000100,
    32'b11001011001110001010001101101001,
    32'b11001010111100010010011001001111,
    32'b11001010101010011010100100110100,
    32'b11001010011000100010110000011010,
    32'b11001010000110101010111011111111,
    32'b11001001110100110011000111100100,
    32'b11001001100010111011010011001010,
    32'b11001001010001000011011110101111,
    32'b11001000111111001011101010010101,
    32'b11001000101101010011110101111010,
    32'b11001000011011011100000001100000,
    32'b11001000001001100100001101000101,
    32'b11000111110111101100011000101011,
    32'b11000111100101110100100100010000,
    32'b11000111010011111100101111110110,
    32'b11000111000010000100111011011011,
    32'b11000110110000001101000111000001,
    32'b11000110011110010101010010100110,
    32'b11000110001100011101011110001011,
    32'b11000101111010100101101001110001,
    32'b11000101101000101101110101010110,
    32'b11000101010110110110000000111100,
    32'b11000101000100111110001100100001,
    32'b11000100110011000110011000000111,
    32'b11000100100001001110100011101100,
    32'b11000100001111010110101111010010,
    32'b11000011111101011110111010110111,
    32'b11000011101011100111000110011101,
    32'b11000011011001101111010010000010,
    32'b11000011000111110111011101101000,
    32'b11000010110101111111101001001101,
    32'b11000010100100000111110100110011,
    32'b11000010010010010000000000011000,
    32'b11000010000000011000001011111101,
    32'b11000001101110100000010111100011,
    32'b11000001011100101000100011001000,
    32'b11000001001010110000101110101110,
    32'b11000000111000111000111010010011,
    32'b11000000100111000001000101111001,
    32'b11000000010101001001010001011110,
    32'b11000000000011010001011101000100,
    32'b10111111110001011001101000101001,
    32'b10111111011111100001110100001111,
    32'b10111111001101101001111111110100,
    32'b10111110111011110010001011011010,
    32'b10111110101001111010010110111111,
    32'b10111110011000000010100010100100,
    32'b10111110000110001010101110001010,
    32'b10111101110100010010111001101111,
    32'b10111101100010011011000101010101,
    32'b10111101010000100011010000111010,
    32'b10111100111110101011011100100000,
    32'b10111100101100110011101000000101,
    32'b10111100011010111011110011101011,
    32'b10111100001001000011111111010000,
    32'b10111011110111001100001010110110,
    32'b10111011100101010100010110011011,
    32'b10111011010011011100100010000001,
    32'b10111011000001100100101101100110,
    32'b10111010101111101100111001001011,
    32'b10111010011101110101000100110001,
    32'b10111010001011111101010000010110,
    32'b10111001111010000101011011111100,
    32'b10111001101000001101100111100001,
    32'b10111001010110010101110011000111,
    32'b10111001000100011101111110101100,
    32'b10111000110010100110001010010010,
    32'b10111000100000101110010101110111,
    32'b10111000001110110110100001011101,
    32'b10110111111100111110101101000010,
    32'b10110111101011000110111000101000,
    32'b10110111011001001111000100001101,
    32'b10110111000111010111001111110011,
    32'b10110110110101011111011011011000,
    32'b10110110100011100111100110111101,
    32'b10110110010001101111110010100011,
    32'b10110101111111110111111110001000,
    32'b10110101101110000000001001101110,
    32'b10110101011100001000010101010011,
    32'b10110101001010010000100000111001,
    32'b10110100111000011000101100011110,
    32'b10110100100110100000111000000100,
    32'b10110100010100101001000011101001,
    32'b10110100000010110001001111001111,
    32'b10110011110000111001011010110100,
    32'b10110011011111000001100110011010,
    32'b10110011001101001001110001111111,
    32'b10110010111011010001111101100100,
    32'b10110010101001011010001001001010,
    32'b10110010010111100010010100101111,
    32'b10110010000101101010100000010101,
    32'b10110001110011110010101011111010,
    32'b10110001100001111010110111100000,
    32'b10110001010000000011000011000101,
    32'b10110000111110001011001110101011,
    32'b10110000101100010011011010010000,
    32'b10110000011010011011100101110110,
    32'b10110000001000100011110001011011,
    32'b10101111110110101011111101000001,
    32'b10101111100100110100001000100110,
    32'b10101111010010111100010100001100,
    32'b10101111000001000100011111110001,
    32'b10101110101111001100101011010110,
    32'b10101110011101010100110110111100,
    32'b10101110001011011101000010100001,
    32'b10101101111001100101001110000111,
    32'b10101101100111101101011001101100,
    32'b10101101010101110101100101010010,
    32'b10101101000011111101110000110111,
    32'b10101100110010000101111100011101,
    32'b10101100100000001110001000000010,
    32'b10101100001110010110010011101000,
    32'b10101011111100011110011111001101,
    32'b10101011101010100110101010110011,
    32'b10101011011000101110110110011000,
    32'b10101011000110110111000001111101,
    32'b10101010110100111111001101100011,
    32'b10101010100011000111011001001000,
    32'b10101010010001001111100100101110,
    32'b10101001111111010111110000010011,
    32'b10101001101101011111111011111001,
    32'b10101001011011101000000111011110,
    32'b10101001001001110000010011000100,
    32'b10101000110111111000011110101001,
    32'b10101000100110000000101010001111,
    32'b10101000010100001000110101110100,
    32'b10101000000010010001000001011010,
    32'b10100111110000011001001100111111,
    32'b10100111011110100001011000100100,
    32'b10100111001100101001100100001010,
    32'b10100110111010110001101111101111,
    32'b10100110101000111001111011010101,
    32'b10100110010111000010000110111010,
    32'b10100110000101001010010010100000,
    32'b10100101110011010010011110000101,
    32'b10100101100001011010101001101011,
    32'b10100101001111100010110101010000,
    32'b10100100111101101011000000110110,
    32'b10100100101011110011001100011011,
    32'b10100100011001111011011000000001,
    32'b10100100001000000011100011100110,
    32'b10100011110110001011101111001100,
    32'b10100011100100010011111010110001,
    32'b10100011010010011100000110010110,
    32'b10100011000000100100010001111100,
    32'b10100010101110101100011101100001,
    32'b10100010011100110100101001000111,
    32'b10100010001010111100110100101100,
    32'b10100001111001000101000000010010,
    32'b10100001100111001101001011110111,
    32'b10100001010101010101010111011101,
    32'b10100001000011011101100011000010,
    32'b10100000110001100101101110101000,
    32'b10100000011111101101111010001101,
    32'b10100000001101110110000101110011,
    32'b10011111111011111110010001011000,
    32'b10011111101010000110011100111101,
    32'b10011111011000001110101000100011,
    32'b10011111000110010110110100001000,
    32'b10011110110100011110111111101110,
    32'b10011110100010100111001011010011,
    32'b10011110010000101111010110111001,
    32'b10011101111110110111100010011110,
    32'b10011101101100111111101110000100,
    32'b10011101011011000111111001101001,
    32'b10011101001001010000000101001111,
    32'b10011100110111011000010000110100,
    32'b10011100100101100000011100011010,
    32'b10011100010011101000100111111111,
    32'b10011100000001110000110011100101,
    32'b10011011101111111000111111001010
  };

  logic [31 : 0] pos_radians [360] = {
    32'b00000000000000000000000000000000,
    32'b00000000010001110111110100011010,
    32'b00000000100011101111101000110101,
    32'b00000000110101100111011101001111,
    32'b00000001000111011111010001101010,
    32'b00000001011001010111000110000100,
    32'b00000001101011001110111010011111,
    32'b00000001111101000110101110111001,
    32'b00000010001110111110100011010100,
    32'b00000010100000110110010111101110,
    32'b00000010110010101110001100001001,
    32'b00000011000100100110000000100011,
    32'b00000011010110011101110100111110,
    32'b00000011101000010101101001011000,
    32'b00000011111010001101011101110011,
    32'b00000100001100000101010010001110,
    32'b00000100011101111101000110101000,
    32'b00000100101111110100111011000011,
    32'b00000101000001101100101111011101,
    32'b00000101010011100100100011111000,
    32'b00000101100101011100011000010010,
    32'b00000101110111010100001100101101,
    32'b00000110001001001100000001000111,
    32'b00000110011011000011110101100010,
    32'b00000110101100111011101001111100,
    32'b00000110111110110011011110010111,
    32'b00000111010000101011010010110001,
    32'b00000111100010100011000111001100,
    32'b00000111110100011010111011100111,
    32'b00001000000110010010110000000001,
    32'b00001000011000001010100100011100,
    32'b00001000101010000010011000110110,
    32'b00001000111011111010001101010001,
    32'b00001001001101110010000001101011,
    32'b00001001011111101001110110000110,
    32'b00001001110001100001101010100000,
    32'b00001010000011011001011110111011,
    32'b00001010010101010001010011010101,
    32'b00001010100111001001000111110000,
    32'b00001010111001000000111100001010,
    32'b00001011001010111000110000100101,
    32'b00001011011100110000100100111111,
    32'b00001011101110101000011001011010,
    32'b00001100000000100000001101110101,
    32'b00001100010010011000000010001111,
    32'b00001100100100001111110110101010,
    32'b00001100110110000111101011000100,
    32'b00001101000111111111011111011111,
    32'b00001101011001110111010011111001,
    32'b00001101101011101111001000010100,
    32'b00001101111101100110111100101110,
    32'b00001110001111011110110001001001,
    32'b00001110100001010110100101100011,
    32'b00001110110011001110011001111110,
    32'b00001111000101000110001110011000,
    32'b00001111010110111110000010110011,
    32'b00001111101000110101110111001110,
    32'b00001111111010101101101011101000,
    32'b00010000001100100101100000000011,
    32'b00010000011110011101010100011101,
    32'b00010000110000010101001000111000,
    32'b00010001000010001100111101010010,
    32'b00010001010100000100110001101101,
    32'b00010001100101111100100110000111,
    32'b00010001110111110100011010100010,
    32'b00010010001001101100001110111100,
    32'b00010010011011100100000011010111,
    32'b00010010101101011011110111110001,
    32'b00010010111111010011101100001100,
    32'b00010011010001001011100000100111,
    32'b00010011100011000011010101000001,
    32'b00010011110100111011001001011100,
    32'b00010100000110110010111101110110,
    32'b00010100011000101010110010010001,
    32'b00010100101010100010100110101011,
    32'b00010100111100011010011011000110,
    32'b00010101001110010010001111100000,
    32'b00010101100000001010000011111011,
    32'b00010101110010000001111000010101,
    32'b00010110000011111001101100110000,
    32'b00010110010101110001100001001010,
    32'b00010110100111101001010101100101,
    32'b00010110111001100001001001111111,
    32'b00010111001011011000111110011010,
    32'b00010111011101010000110010110101,
    32'b00010111101111001000100111001111,
    32'b00011000000001000000011011101010,
    32'b00011000010010111000010000000100,
    32'b00011000100100110000000100011111,
    32'b00011000110110100111111000111001,
    32'b00011001001000011111101101010100,
    32'b00011001011010010111100001101110,
    32'b00011001101100001111010110001001,
    32'b00011001111110000111001010100011,
    32'b00011010001111111110111110111110,
    32'b00011010100001110110110011011000,
    32'b00011010110011101110100111110011,
    32'b00011011000101100110011100001110,
    32'b00011011010111011110010000101000,
    32'b00011011101001010110000101000011,
    32'b00011011111011001101111001011101,
    32'b00011100001101000101101101111000,
    32'b00011100011110111101100010010010,
    32'b00011100110000110101010110101101,
    32'b00011101000010101101001011000111,
    32'b00011101010100100100111111100010,
    32'b00011101100110011100110011111100,
    32'b00011101111000010100101000010111,
    32'b00011110001010001100011100110001,
    32'b00011110011100000100010001001100,
    32'b00011110101101111100000101100110,
    32'b00011110111111110011111010000001,
    32'b00011111010001101011101110011100,
    32'b00011111100011100011100010110110,
    32'b00011111110101011011010111010001,
    32'b00100000000111010011001011101011,
    32'b00100000011001001011000000000110,
    32'b00100000101011000010110100100000,
    32'b00100000111100111010101000111011,
    32'b00100001001110110010011101010101,
    32'b00100001100000101010010001110000,
    32'b00100001110010100010000110001010,
    32'b00100010000100011001111010100101,
    32'b00100010010110010001101110111111,
    32'b00100010101000001001100011011010,
    32'b00100010111010000001010111110101,
    32'b00100011001011111001001100001111,
    32'b00100011011101110001000000101010,
    32'b00100011101111101000110101000100,
    32'b00100100000001100000101001011111,
    32'b00100100010011011000011101111001,
    32'b00100100100101010000010010010100,
    32'b00100100110111001000000110101110,
    32'b00100101001000111111111011001001,
    32'b00100101011010110111101111100011,
    32'b00100101101100101111100011111110,
    32'b00100101111110100111011000011000,
    32'b00100110010000011111001100110011,
    32'b00100110100010010111000001001110,
    32'b00100110110100001110110101101000,
    32'b00100111000110000110101010000011,
    32'b00100111010111111110011110011101,
    32'b00100111101001110110010010111000,
    32'b00100111111011101110000111010010,
    32'b00101000001101100101111011101101,
    32'b00101000011111011101110000000111,
    32'b00101000110001010101100100100010,
    32'b00101001000011001101011000111100,
    32'b00101001010101000101001101010111,
    32'b00101001100110111101000001110001,
    32'b00101001111000110100110110001100,
    32'b00101010001010101100101010100110,
    32'b00101010011100100100011111000001,
    32'b00101010101110011100010011011100,
    32'b00101011000000010100000111110110,
    32'b00101011010010001011111100010001,
    32'b00101011100100000011110000101011,
    32'b00101011110101111011100101000110,
    32'b00101100000111110011011001100000,
    32'b00101100011001101011001101111011,
    32'b00101100101011100011000010010101,
    32'b00101100111101011010110110110000,
    32'b00101101001111010010101011001010,
    32'b00101101100001001010011111100101,
    32'b00101101110011000010010011111111,
    32'b00101110000100111010001000011010,
    32'b00101110010110110001111100110101,
    32'b00101110101000101001110001001111,
    32'b00101110111010100001100101101010,
    32'b00101111001100011001011010000100,
    32'b00101111011110010001001110011111,
    32'b00101111110000001001000010111001,
    32'b00110000000010000000110111010100,
    32'b00110000010011111000101011101110,
    32'b00110000100101110000100000001001,
    32'b00110000110111101000010100100011,
    32'b00110001001001100000001000111110,
    32'b00110001011011010111111101011000,
    32'b00110001101101001111110001110011,
    32'b00110001111111000111100110001101,
    32'b00110010010000111111011010101000,
    32'b00110010100010110111001111000011,
    32'b00110010110100101111000011011101,
    32'b00110011000110100110110111111000,
    32'b00110011011000011110101100010010,
    32'b00110011101010010110100000101101,
    32'b00110011111100001110010101000111,
    32'b00110100001110000110001001100010,
    32'b00110100011111111101111101111100,
    32'b00110100110001110101110010010111,
    32'b00110101000011101101100110110001,
    32'b00110101010101100101011011001100,
    32'b00110101100111011101001111100110,
    32'b00110101111001010101000100000001,
    32'b00110110001011001100111000011100,
    32'b00110110011101000100101100110110,
    32'b00110110101110111100100001010001,
    32'b00110111000000110100010101101011,
    32'b00110111010010101100001010000110,
    32'b00110111100100100011111110100000,
    32'b00110111110110011011110010111011,
    32'b00111000001000010011100111010101,
    32'b00111000011010001011011011110000,
    32'b00111000101100000011010000001010,
    32'b00111000111101111011000100100101,
    32'b00111001001111110010111000111111,
    32'b00111001100001101010101101011010,
    32'b00111001110011100010100001110101,
    32'b00111010000101011010010110001111,
    32'b00111010010111010010001010101010,
    32'b00111010101001001001111111000100,
    32'b00111010111011000001110011011111,
    32'b00111011001100111001100111111001,
    32'b00111011011110110001011100010100,
    32'b00111011110000101001010000101110,
    32'b00111100000010100001000101001001,
    32'b00111100010100011000111001100011,
    32'b00111100100110010000101101111110,
    32'b00111100111000001000100010011000,
    32'b00111101001010000000010110110011,
    32'b00111101011011111000001011001101,
    32'b00111101101101101111111111101000,
    32'b00111101111111100111110100000011,
    32'b00111110010001011111101000011101,
    32'b00111110100011010111011100111000,
    32'b00111110110101001111010001010010,
    32'b00111111000111000111000101101101,
    32'b00111111011000111110111010000111,
    32'b00111111101010110110101110100010,
    32'b00111111111100101110100010111100,
    32'b01000000001110100110010111010111,
    32'b01000000100000011110001011110001,
    32'b01000000110010010110000000001100,
    32'b01000001000100001101110100100110,
    32'b01000001010110000101101001000001,
    32'b01000001100111111101011101011100,
    32'b01000001111001110101010001110110,
    32'b01000010001011101101000110010001,
    32'b01000010011101100100111010101011,
    32'b01000010101111011100101111000110,
    32'b01000011000001010100100011100000,
    32'b01000011010011001100010111111011,
    32'b01000011100101000100001100010101,
    32'b01000011110110111100000000110000,
    32'b01000100001000110011110101001010,
    32'b01000100011010101011101001100101,
    32'b01000100101100100011011101111111,
    32'b01000100111110011011010010011010,
    32'b01000101010000010011000110110101,
    32'b01000101100010001010111011001111,
    32'b01000101110100000010101111101010,
    32'b01000110000101111010100100000100,
    32'b01000110010111110010011000011111,
    32'b01000110101001101010001100111001,
    32'b01000110111011100010000001010100,
    32'b01000111001101011001110101101110,
    32'b01000111011111010001101010001001,
    32'b01000111110001001001011110100011,
    32'b01001000000011000001010010111110,
    32'b01001000010100111001000111011000,
    32'b01001000100110110000111011110011,
    32'b01001000111000101000110000001101,
    32'b01001001001010100000100100101000,
    32'b01001001011100011000011001000011,
    32'b01001001101110010000001101011101,
    32'b01001010000000001000000001111000,
    32'b01001010010001111111110110010010,
    32'b01001010100011110111101010101101,
    32'b01001010110101101111011111000111,
    32'b01001011000111100111010011100010,
    32'b01001011011001011111000111111100,
    32'b01001011101011010110111100010111,
    32'b01001011111101001110110000110001,
    32'b01001100001111000110100101001100,
    32'b01001100100000111110011001100110,
    32'b01001100110010110110001110000001,
    32'b01001101000100101110000010011100,
    32'b01001101010110100101110110110110,
    32'b01001101101000011101101011010001,
    32'b01001101111010010101011111101011,
    32'b01001110001100001101010100000110,
    32'b01001110011110000101001000100000,
    32'b01001110101111111100111100111011,
    32'b01001111000001110100110001010101,
    32'b01001111010011101100100101110000,
    32'b01001111100101100100011010001010,
    32'b01001111110111011100001110100101,
    32'b01010000001001010100000010111111,
    32'b01010000011011001011110111011010,
    32'b01010000101101000011101011110100,
    32'b01010000111110111011100000001111,
    32'b01010001010000110011010100101010,
    32'b01010001100010101011001001000100,
    32'b01010001110100100010111101011111,
    32'b01010010000110011010110001111001,
    32'b01010010011000010010100110010100,
    32'b01010010101010001010011010101110,
    32'b01010010111100000010001111001001,
    32'b01010011001101111010000011100011,
    32'b01010011011111110001110111111110,
    32'b01010011110001101001101100011000,
    32'b01010100000011100001100000110011,
    32'b01010100010101011001010101001101,
    32'b01010100100111010001001001101000,
    32'b01010100111001001000111110000011,
    32'b01010101001011000000110010011101,
    32'b01010101011100111000100110111000,
    32'b01010101101110110000011011010010,
    32'b01010110000000101000001111101101,
    32'b01010110010010100000000100000111,
    32'b01010110100100010111111000100010,
    32'b01010110110110001111101100111100,
    32'b01010111001000000111100001010111,
    32'b01010111011001111111010101110001,
    32'b01010111101011110111001010001100,
    32'b01010111111101101110111110100110,
    32'b01011000001111100110110011000001,
    32'b01011000100001011110100111011100,
    32'b01011000110011010110011011110110,
    32'b01011001000101001110010000010001,
    32'b01011001010111000110000100101011,
    32'b01011001101000111101111001000110,
    32'b01011001111010110101101101100000,
    32'b01011010001100101101100001111011,
    32'b01011010011110100101010110010101,
    32'b01011010110000011101001010110000,
    32'b01011011000010010100111111001010,
    32'b01011011010100001100110011100101,
    32'b01011011100110000100100111111111,
    32'b01011011110111111100011100011010,
    32'b01011100001001110100010000110100,
    32'b01011100011011101100000101001111,
    32'b01011100101101100011111001101010,
    32'b01011100111111011011101110000100,
    32'b01011101010001010011100010011111,
    32'b01011101100011001011010110111001,
    32'b01011101110101000011001011010100,
    32'b01011110000110111010111111101110,
    32'b01011110011000110010110100001001,
    32'b01011110101010101010101000100011,
    32'b01011110111100100010011100111110,
    32'b01011111001110011010010001011000,
    32'b01011111100000010010000101110011,
    32'b01011111110010001001111010001101,
    32'b01100000000100000001101110101000,
    32'b01100000010101111001100011000011,
    32'b01100000100111110001010111011101,
    32'b01100000111001101001001011111000,
    32'b01100001001011100001000000010010,
    32'b01100001011101011000110100101101,
    32'b01100001101111010000101001000111,
    32'b01100010000001001000011101100010,
    32'b01100010010011000000010001111100,
    32'b01100010100100111000000110010111,
    32'b01100010110110101111111010110001,
    32'b01100011001000100111101111001100,
    32'b01100011011010011111100011100110,
    32'b01100011101100010111011000000001,
    32'b01100011111110001111001100011011,
    32'b01100100010000000111000000110110
  };

endpackage

`endif
