import vip_axi4s_types_pkg::*;

`include "vip_axi4s_pkg.sv"
`include "vip_axi4s_if.sv"
