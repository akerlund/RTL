module dummy();
endmodule