////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2020 Fredrik Åkerlund
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <https://www.gnu.org/licenses/>.
//
// Description:
//
////////////////////////////////////////////////////////////////////////////////

class clk_rst_item extends uvm_sequence_item;

  reset_edge_t  reset_edge  = RESET_AT_CLK_RISING_EDGE_E;
  reset_value_t reset_value = RESET_INACTIVE_E;

  `uvm_object_utils(clk_rst_item)

  function new(string name = "clk_rst_item");
    super.new(name);
  endfunction

endclass
