package gf_ref_pkg;

localparam int M_C        = 8;
localparam int P_ORDER_C  = 256;
localparam int REF_SIZE_C = 16;

localparam logic [M_C-1 : 0] GF_ADD_C [REF_SIZE_C] [3] = '{
  '{158,150,8},
  '{208,16,192},
  '{96,25,121},
  '{36,163,135},
  '{121,230,159},
  '{252,33,221},
  '{47,24,55},
  '{17,14,31},
  '{92,204,144},
  '{234,77,167},
  '{21,75,94},
  '{24,76,84},
  '{1,212,213},
  '{220,2,222},
  '{59,140,183},
  '{189,55,138}
};

localparam logic [M_C-1 : 0] GF_MUL_C [REF_SIZE_C] [3] = '{
  '{147,26,58},
  '{81,204,115},
  '{57,65,251},
  '{213,137,158},
  '{236,221,39},
  '{101,31,47},
  '{54,3,90},
  '{3,133,148},
  '{88,104,242},
  '{149,209,136},
  '{227,31,116},
  '{42,170,244},
  '{212,132,68},
  '{127,171,210},
  '{96,157,106},
  '{69,87,12}
};

localparam logic [M_C-1 : 0] GF_DIV_C [REF_SIZE_C] [3] = '{
  '{8,46,103},
  '{136,248,103},
  '{0,105,0},
  '{229,79,140},
  '{214,48,26},
  '{156,126,132},
  '{132,76,232},
  '{46,253,225},
  '{105,244,239},
  '{181,228,110},
  '{103,163,74},
  '{198,191,205},
  '{64,3,201},
  '{97,147,124},
  '{171,16,27},
  '{211,19,230}
};

endpackage
